
module fsmir (
	input              clk   ,
	input        [7:0] di    ,
	output logic [7:0] c     ,
	output             solved
);

	initial c = 8'b0;

	assign solved = c == 8'd59;

	always @(posedge clk) begin
		c <= 8'b0;

		case (c)

			8'b1001: if((di ^ c) == 8'b1110000) c <= 8'b1010;
			8'b101001: if((di ^ c) == 8'b1010000) c <= 8'b101010;
			8'b11100: if((di ^ c) == 8'b1101000) c <= 8'b11101;
			8'b1010: if((di ^ c) == 8'b1111001) c <= 8'b1011;
			8'b1100: if((di ^ c) == 8'b1101001) c <= 8'b1101;
			8'b110000: if((di ^ c) == 8'b1011001) c <= 8'b110001;
			8'b111001: if((di ^ c) == 8'b110) c <= 8'b111010;
			8'b11000: if((di ^ c) == 8'b1000111) c <= 8'b11001;
			8'b11110: if((di ^ c) == 8'b1011101) c <= 8'b11111;
			8'b10: if((di ^ c) == 8'b1110001) c <= 8'b11;
			8'b10100: if((di ^ c) == 8'b1110011) c <= 8'b10101;
			8'b101011: if((di ^ c) == 8'b1000101) c <= 8'b101100;
			8'b10000: if((di ^ c) == 8'b1100010) c <= 8'b10001;
			8'b101010: if((di ^ c) == 8'b1110101) c <= 8'b101011;
			8'b100111: if((di ^ c) == 8'b1001001) c <= 8'b101000;
			8'b10111: if((di ^ c) == 8'b1100100) c <= 8'b11000;
			8'b11: if((di ^ c) == 8'b1110111) c <= 8'b100;
			8'b1111: if((di ^ c) == 8'b1101010) c <= 8'b10000;
			8'b101101: if((di ^ c) == 8'b1011001) c <= 8'b101110;
			8'b101000: if((di ^ c) == 8'b1001011) c <= 8'b101001;
			8'b101: if((di ^ c) == 8'b1010001) c <= 8'b110;
			8'b110110: if((di ^ c) == 8'b1010001) c <= 8'b110111;
			8'b1110: if((di ^ c) == 8'b1011000) c <= 8'b1111;
			8'b100010: if((di ^ c) == 8'b1010110) c <= 8'b100011;
			8'b100101: if((di ^ c) == 8'b1000011) c <= 8'b100110;
			8'b100: if((di ^ c) == 8'b1000111) c <= 8'b101;
			8'b10010: if((di ^ c) == 8'b1111110) c <= 8'b10011;
			8'b1101: if((di ^ c) == 8'b1100000) c <= 8'b1110;
			8'b110001: if((di ^ c) == 8'b1011110) c <= 8'b110010;
			8'b110101: if((di ^ c) == 8'b1011100) c <= 8'b110110;
			8'b110011: if((di ^ c) == 8'b1101100) c <= 8'b110100;
			8'b101111: if((di ^ c) == 8'b1011011) c <= 8'b110000;
			8'b1: if((di ^ c) == 8'b1110100) c <= 8'b10;
			8'b11001: if((di ^ c) == 8'b1110011) c <= 8'b11010;
			8'b100000: if((di ^ c) == 8'b1010111) c <= 8'b100001;
			8'b100011: if((di ^ c) == 8'b1001011) c <= 8'b100100;
			8'b100100: if((di ^ c) == 8'b1111011) c <= 8'b100101;
			8'b110111: if((di ^ c) == 8'b1011111) c <= 8'b111000;
			8'b100001: if((di ^ c) == 8'b1001000) c <= 8'b100010;
			8'b11101: if((di ^ c) == 8'b1000010) c <= 8'b11110;
			8'b110: if((di ^ c) == 8'b1000000) c <= 8'b111;
			8'b1000: if((di ^ c) == 8'b1011011) c <= 8'b1001;
			8'b110010: if((di ^ c) == 8'b1011100) c <= 8'b110011;
			8'b10011: if((di ^ c) == 8'b1111100) c <= 8'b10100;
			8'b100110: if((di ^ c) == 8'b1000111) c <= 8'b100111;
			8'b111010: if((di ^ c) == 8'b1000111) c <= 8'b111011;
			8'b10001: if((di ^ c) == 8'b1111000) c <= 8'b10010;
			8'b10101: if((di ^ c) == 8'b1001010) c <= 8'b10110;
			8'b0: if((di ^ c) == 8'b1101010) c <= 8'b1;
			8'b111000: if((di ^ c) == 8'b1001100) c <= 8'b111001;
			8'b110100: if((di ^ c) == 8'b1000110) c <= 8'b110101;
			8'b1011: if((di ^ c) == 8'b1111111) c <= 8'b1100;
			8'b11011: if((di ^ c) == 8'b1101000) c <= 8'b11100;
			8'b11111: if((di ^ c) == 8'b1000000) c <= 8'b100000;
			8'b101110: if((di ^ c) == 8'b1001111) c <= 8'b101111;
			8'b10110: if((di ^ c) == 8'b1111111) c <= 8'b10111;
			8'b11010: if((di ^ c) == 8'b1101111) c <= 8'b11011;
			8'b111: if((di ^ c) == 8'b1111100) c <= 8'b1000;
			8'b101100: if((di ^ c) == 8'b1000011) c <= 8'b101101;

			default   : c <= 8'b0;
		endcase
	end
endmodule

