	assign solved = c == 9'b101001101;
			9'b0 : case(di)
				8'b1000011: c <= 9'b1011010;
				8'b101000: c <= 9'b10111010;
				8'b111010: c <= 9'b100000110;
				8'b110110: c <= 9'b110010011;
				8'b1100100: c <= 9'b111010110;
				8'b1000000: c <= 9'b101000100;
				8'b1110110: c <= 9'b101011;
				8'b100101: c <= 9'b11001110;
				8'b101111: c <= 9'b100000011;
				8'b100110: c <= 9'b11101111;
				8'b1100011: c <= 9'b100110100;
				8'b1001000: c <= 9'b100000010;
				8'b111000: c <= 9'b111011;
				8'b110001: c <= 9'b100001001;
				8'b1010111: c <= 9'b11111110;
				8'b1001110: c <= 9'b10101;
				8'b1101010: c <= 9'b111110010;
				8'b1001001: c <= 9'b11100111;
				8'b1100000: c <= 9'b1100001;
				8'b110111: c <= 9'b100000111;
				8'b1011101: c <= 9'b100110010;
				8'b1011011: c <= 9'b11000;
				8'b111001: c <= 9'b111101010;
				8'b1001010: c <= 9'b111;
				8'b110011: c <= 9'b11010100;
				8'b1101100: c <= 9'b11001000;
				8'b1110111: c <= 9'b101101111;
				8'b101011: c <= 9'b10100;
				8'b1101011: c <= 9'b10101101;
				8'b111100: c <= 9'b10001000;
				8'b1000111: c <= 9'b111111110;
				8'b1011111: c <= 9'b111001110;
				8'b1110100: c <= 9'b10101000;
				8'b101101: c <= 9'b111010110;
				8'b1010011: c <= 9'b101110010;
				8'b1100001: c <= 9'b10110010;
				8'b110101: c <= 9'b110100010;
				8'b1000100: c <= 9'b101001000;
				8'b1010001: c <= 9'b101101100;
				8'b1010100: c <= 9'b10001011;
				8'b1100110: c <= 9'b101101010;
				8'b101010: c <= 9'b11100101;
				8'b1011110: c <= 9'b110110011;
				8'b1100111: c <= 9'b11000011;
				8'b1011010: c <= 9'b111101001;
				8'b1000010: c <= 9'b101011000;
				8'b111101: c <= 9'b1011000;
				8'b110000: c <= 9'b111111110;
				8'b111110: c <= 9'b110001011;
				8'b1100010: c <= 9'b101100000;
				8'b1110000: c <= 9'b100000101;
				8'b1101001: c <= 9'b110101101;
				8'b1110011: c <= 9'b100001011;
				8'b1001100: c <= 9'b110101001;
				8'b100001: c <= 9'b101000010;
				8'b1000110: c <= 9'b101001000;
				8'b1110010: c <= 9'b111011;
				8'b1010000: c <= 9'b1000010;
				8'b1111010: c <= 9'b100100000;
				8'b1010101: c <= 9'b110;
				8'b111011: c <= 9'b101010011;
				8'b1001101: c <= 9'b1110001;
				8'b111111: c <= 9'b111111110;
				8'b1101110: c <= 9'b100101101;
				8'b1111011: c <= 9'b1110100;
				8'b1001011: c <= 9'b110111000;
				8'b1101111: c <= 9'b100110010;
				8'b1101000: c <= 9'b100000010;
				8'b101100: c <= 9'b101010111;
				8'b100100: c <= 9'b100010010;
				8'b1111000: c <= 9'b101;
				8'b1000101: c <= 9'b1110100;
				8'b1011001: c <= 9'b110;
				8'b110100: c <= 9'b10110011;
				8'b1111001: c <= 9'b110111;
				8'b1110001: c <= 9'b1100010;
				8'b1001111: c <= 9'b11110110;
				8'b1100101: c <= 9'b100010110;
				8'b1111110: c <= 9'b101100010;
				8'b1111100: c <= 9'b100110111;
				8'b1010110: c <= 9'b1110000;
				8'b110010: c <= 9'b110100000;
				8'b1101101: c <= 9'b111011011;
				8'b100011: c <= 9'b101001111;
				8'b1110101: c <= 9'b110100101;
				8'b1111101: c <= 9'b10001000;
				8'b101001: c <= 9'b10111110;
				8'b1010010: c <= 9'b11;
				8'b1011000: c <= 9'b100101010;
				8'b101110: c <= 9'b10001100;
				8'b1000001: c <= 9'b11001011;
				default: c <= 9'b0;
			endcase
			9'b111110010 : case(di)
				8'b1000011: c <= 9'b100110011;
				8'b101000: c <= 9'b100000111;
				8'b111010: c <= 9'b110011111;
				8'b110110: c <= 9'b101100000;
				8'b1100100: c <= 9'b100101010;
				8'b1000000: c <= 9'b10001110;
				8'b1110110: c <= 9'b111111;
				8'b100101: c <= 9'b1001001;
				8'b101111: c <= 9'b111101010;
				8'b100110: c <= 9'b11100010;
				8'b1100011: c <= 9'b111100111;
				8'b1001000: c <= 9'b11001000;
				8'b111000: c <= 9'b11100011;
				8'b110001: c <= 9'b101110;
				8'b1010111: c <= 9'b10101001;
				8'b1001110: c <= 9'b110001111;
				8'b1101010: c <= 9'b10000111;
				8'b1001001: c <= 9'b11001111;
				8'b1100000: c <= 9'b11001100;
				8'b110111: c <= 9'b10110001;
				8'b1011101: c <= 9'b100000101;
				8'b1011011: c <= 9'b111100111;
				8'b111001: c <= 9'b1111111;
				8'b1001010: c <= 9'b10011001;
				8'b110011: c <= 9'b110000110;
				8'b1101100: c <= 9'b11000010;
				8'b1110111: c <= 9'b100010011;
				8'b101011: c <= 9'b100010101;
				8'b1101011: c <= 9'b10110010;
				8'b111100: c <= 9'b10100010;
				8'b1000111: c <= 9'b11000100;
				8'b1011111: c <= 9'b110011011;
				8'b1110100: c <= 9'b111100111;
				8'b101101: c <= 9'b110000001;
				8'b1010011: c <= 9'b111101111;
				8'b1100001: c <= 9'b101110100;
				8'b110101: c <= 9'b1111001;
				8'b1000100: c <= 9'b1001001;
				8'b1010001: c <= 9'b1000001;
				8'b1010100: c <= 9'b110100101;
				8'b1100110: c <= 9'b101000011;
				8'b101010: c <= 9'b101110101;
				8'b1011110: c <= 9'b10101010;
				8'b1100111: c <= 9'b101010010;
				8'b1011010: c <= 9'b100011111;
				8'b1000010: c <= 9'b1011100;
				8'b111101: c <= 9'b111011101;
				8'b110000: c <= 9'b1010111;
				8'b111110: c <= 9'b101100010;
				8'b1100010: c <= 9'b1110100;
				8'b1110000: c <= 9'b10010;
				8'b1101001: c <= 9'b100110110;
				8'b1110011: c <= 9'b110111010;
				8'b1001100: c <= 9'b110000000;
				8'b100001: c <= 9'b100000010;
				8'b1000110: c <= 9'b110011101;
				8'b1110010: c <= 9'b100101110;
				8'b1010000: c <= 9'b1111111;
				8'b1111010: c <= 9'b100101001;
				8'b1010101: c <= 9'b101000100;
				8'b111011: c <= 9'b1011001;
				8'b1001101: c <= 9'b11000010;
				8'b111111: c <= 9'b1010010;
				8'b1101110: c <= 9'b1011011;
				8'b1111011: c <= 9'b11011100;
				8'b1001011: c <= 9'b101001100;
				8'b1101111: c <= 9'b110011001;
				8'b1101000: c <= 9'b101111110;
				8'b101100: c <= 9'b110101100;
				8'b100100: c <= 9'b100010;
				8'b1111000: c <= 9'b10001000;
				8'b1000101: c <= 9'b110100100;
				8'b1011001: c <= 9'b10100111;
				8'b110100: c <= 9'b1101110;
				8'b1111001: c <= 9'b10100111;
				8'b1110001: c <= 9'b1010011;
				8'b1001111: c <= 9'b1010101;
				8'b1100101: c <= 9'b1111110;
				8'b1111110: c <= 9'b101001100;
				8'b1111100: c <= 9'b1100;
				8'b1010110: c <= 9'b111110011;
				8'b110010: c <= 9'b1111101;
				8'b1101101: c <= 9'b100100001;
				8'b100011: c <= 9'b101010111;
				8'b1110101: c <= 9'b110101000;
				8'b1111101: c <= 9'b100100110;
				8'b101001: c <= 9'b11;
				8'b1010010: c <= 9'b110100;
				8'b1011000: c <= 9'b11111110;
				8'b101110: c <= 9'b1010001;
				8'b1000001: c <= 9'b11011;
				default: c <= 9'b0;
			endcase
			9'b110101000 : case(di)
				8'b1000011: c <= 9'b10110001;
				8'b101000: c <= 9'b100100;
				8'b111010: c <= 9'b1010000;
				8'b110110: c <= 9'b10100;
				8'b1100100: c <= 9'b11011100;
				8'b1000000: c <= 9'b100010110;
				8'b1110110: c <= 9'b11010001;
				8'b100101: c <= 9'b1000111;
				8'b101111: c <= 9'b10111010;
				8'b100110: c <= 9'b110001101;
				8'b1100011: c <= 9'b100011001;
				8'b1001000: c <= 9'b11110111;
				8'b111000: c <= 9'b1100;
				8'b110001: c <= 9'b110111011;
				8'b1010111: c <= 9'b1010110;
				8'b1001110: c <= 9'b100010011;
				8'b1101010: c <= 9'b111010001;
				8'b1001001: c <= 9'b1100001;
				8'b1100000: c <= 9'b10000001;
				8'b110111: c <= 9'b1000011;
				8'b1011101: c <= 9'b11111000;
				8'b1011011: c <= 9'b1101100;
				8'b111001: c <= 9'b11001100;
				8'b1001010: c <= 9'b11101100;
				8'b110011: c <= 9'b110110010;
				8'b1101100: c <= 9'b1110;
				8'b1110111: c <= 9'b100111010;
				8'b101011: c <= 9'b10001011;
				8'b1101011: c <= 9'b101000010;
				8'b111100: c <= 9'b10111010;
				8'b1000111: c <= 9'b110011;
				8'b1011111: c <= 9'b10111011;
				8'b1110100: c <= 9'b110111001;
				8'b101101: c <= 9'b111101101;
				8'b1010011: c <= 9'b11110001;
				8'b1100001: c <= 9'b10100111;
				8'b110101: c <= 9'b101011001;
				8'b1000100: c <= 9'b11000010;
				8'b1010001: c <= 9'b100;
				8'b1010100: c <= 9'b101110010;
				8'b1100110: c <= 9'b110111110;
				8'b101010: c <= 9'b111010111;
				8'b1011110: c <= 9'b1001100;
				8'b1100111: c <= 9'b100100101;
				8'b1011010: c <= 9'b10001011;
				8'b1000010: c <= 9'b111010111;
				8'b111101: c <= 9'b11111001;
				8'b110000: c <= 9'b101011010;
				8'b111110: c <= 9'b11101100;
				8'b1100010: c <= 9'b100011111;
				8'b1110000: c <= 9'b11110100;
				8'b1101001: c <= 9'b100000111;
				8'b1110011: c <= 9'b100001000;
				8'b1001100: c <= 9'b111011010;
				8'b100001: c <= 9'b11100001;
				8'b1000110: c <= 9'b100110101;
				8'b1110010: c <= 9'b101101000;
				8'b1010000: c <= 9'b110011000;
				8'b1111010: c <= 9'b100111100;
				8'b1010101: c <= 9'b101011;
				8'b111011: c <= 9'b111001010;
				8'b1001101: c <= 9'b110110111;
				8'b111111: c <= 9'b110111110;
				8'b1101110: c <= 9'b111001101;
				8'b1111011: c <= 9'b110000111;
				8'b1001011: c <= 9'b10011011;
				8'b1101111: c <= 9'b11100101;
				8'b1101000: c <= 9'b10011000;
				8'b101100: c <= 9'b100110111;
				8'b100100: c <= 9'b1101010;
				8'b1111000: c <= 9'b101100110;
				8'b1000101: c <= 9'b1001010;
				8'b1011001: c <= 9'b111111111;
				8'b110100: c <= 9'b111001010;
				8'b1111001: c <= 9'b11011110;
				8'b1110001: c <= 9'b11100110;
				8'b1001111: c <= 9'b1111101;
				8'b1100101: c <= 9'b101110001;
				8'b1111110: c <= 9'b100110011;
				8'b1111100: c <= 9'b110010100;
				8'b1010110: c <= 9'b10001001;
				8'b110010: c <= 9'b101011111;
				8'b1101101: c <= 9'b111001101;
				8'b100011: c <= 9'b110101010;
				8'b1110101: c <= 9'b111011110;
				8'b1111101: c <= 9'b100100011;
				8'b101001: c <= 9'b100001010;
				8'b1010010: c <= 9'b110001011;
				8'b1011000: c <= 9'b111101101;
				8'b101110: c <= 9'b11110001;
				8'b1000001: c <= 9'b11111100;
				default: c <= 9'b0;
			endcase
			9'b100001000 : case(di)
				8'b1000011: c <= 9'b10011011;
				8'b101000: c <= 9'b100000110;
				8'b111010: c <= 9'b101100010;
				8'b110110: c <= 9'b11110010;
				8'b1100100: c <= 9'b111110001;
				8'b1000000: c <= 9'b111101010;
				8'b1110110: c <= 9'b111101100;
				8'b100101: c <= 9'b1011110;
				8'b101111: c <= 9'b11100110;
				8'b100110: c <= 9'b100000101;
				8'b1100011: c <= 9'b1011000;
				8'b1001000: c <= 9'b110100110;
				8'b111000: c <= 9'b110001011;
				8'b110001: c <= 9'b100010000;
				8'b1010111: c <= 9'b110110111;
				8'b1001110: c <= 9'b11010111;
				8'b1101010: c <= 9'b100111011;
				8'b1001001: c <= 9'b111100001;
				8'b1100000: c <= 9'b1010010;
				8'b110111: c <= 9'b10110011;
				8'b1011101: c <= 9'b110110;
				8'b1011011: c <= 9'b100101100;
				8'b111001: c <= 9'b1000001;
				8'b1001010: c <= 9'b1111000;
				8'b110011: c <= 9'b1101110;
				8'b1101100: c <= 9'b10111011;
				8'b1110111: c <= 9'b111001001;
				8'b101011: c <= 9'b101001;
				8'b1101011: c <= 9'b10001000;
				8'b111100: c <= 9'b111011;
				8'b1000111: c <= 9'b11101101;
				8'b1011111: c <= 9'b111011100;
				8'b1110100: c <= 9'b110000100;
				8'b101101: c <= 9'b111111010;
				8'b1010011: c <= 9'b10011111;
				8'b1100001: c <= 9'b10111011;
				8'b110101: c <= 9'b10111;
				8'b1000100: c <= 9'b111011111;
				8'b1010001: c <= 9'b111111110;
				8'b1010100: c <= 9'b110000;
				8'b1100110: c <= 9'b11000011;
				8'b101010: c <= 9'b100010011;
				8'b1011110: c <= 9'b11111000;
				8'b1100111: c <= 9'b1010101;
				8'b1011010: c <= 9'b1001110;
				8'b1000010: c <= 9'b1011100;
				8'b111101: c <= 9'b1111000;
				8'b110000: c <= 9'b110001101;
				8'b111110: c <= 9'b1100110;
				8'b1100010: c <= 9'b11111110;
				8'b1110000: c <= 9'b1010101;
				8'b1101001: c <= 9'b11110101;
				8'b1110011: c <= 9'b100000011;
				8'b1001100: c <= 9'b11001011;
				8'b100001: c <= 9'b110001111;
				8'b1000110: c <= 9'b100001101;
				8'b1110010: c <= 9'b11111000;
				8'b1010000: c <= 9'b101010110;
				8'b1111010: c <= 9'b110111111;
				8'b1010101: c <= 9'b11100001;
				8'b111011: c <= 9'b101001;
				8'b1001101: c <= 9'b1011011;
				8'b111111: c <= 9'b1000111;
				8'b1101110: c <= 9'b10001101;
				8'b1111011: c <= 9'b11101011;
				8'b1001011: c <= 9'b111101010;
				8'b1101111: c <= 9'b110000001;
				8'b1101000: c <= 9'b101010010;
				8'b101100: c <= 9'b101111110;
				8'b100100: c <= 9'b11010001;
				8'b1111000: c <= 9'b11110100;
				8'b1000101: c <= 9'b1100100;
				8'b1011001: c <= 9'b1110;
				8'b110100: c <= 9'b110011010;
				8'b1111001: c <= 9'b11001111;
				8'b1110001: c <= 9'b101111111;
				8'b1001111: c <= 9'b10111000;
				8'b1100101: c <= 9'b110100010;
				8'b1111110: c <= 9'b110001110;
				8'b1111100: c <= 9'b1000010;
				8'b1010110: c <= 9'b1101100;
				8'b110010: c <= 9'b10100110;
				8'b1101101: c <= 9'b100000001;
				8'b100011: c <= 9'b1001011;
				8'b1110101: c <= 9'b1001001;
				8'b1111101: c <= 9'b10100100;
				8'b101001: c <= 9'b100111001;
				8'b1010010: c <= 9'b1100100;
				8'b1011000: c <= 9'b11110001;
				8'b101110: c <= 9'b11011110;
				8'b1000001: c <= 9'b100001;
				default: c <= 9'b0;
			endcase
			9'b110000100 : case(di)
				8'b1000011: c <= 9'b1101011;
				8'b101000: c <= 9'b100100;
				8'b111010: c <= 9'b1010111;
				8'b110110: c <= 9'b100100110;
				8'b1100100: c <= 9'b101111000;
				8'b1000000: c <= 9'b10010111;
				8'b1110110: c <= 9'b11100111;
				8'b100101: c <= 9'b111100111;
				8'b101111: c <= 9'b111000;
				8'b100110: c <= 9'b111100001;
				8'b1100011: c <= 9'b10010110;
				8'b1001000: c <= 9'b110010100;
				8'b111000: c <= 9'b111001110;
				8'b110001: c <= 9'b100000010;
				8'b1010111: c <= 9'b100011100;
				8'b1001110: c <= 9'b10011010;
				8'b1101010: c <= 9'b1110010;
				8'b1001001: c <= 9'b1111010;
				8'b1100000: c <= 9'b110000;
				8'b110111: c <= 9'b10011010;
				8'b1011101: c <= 9'b110001111;
				8'b1011011: c <= 9'b11001010;
				8'b111001: c <= 9'b11110101;
				8'b1001010: c <= 9'b10101110;
				8'b110011: c <= 9'b110010010;
				8'b1101100: c <= 9'b10111000;
				8'b1110111: c <= 9'b111011101;
				8'b101011: c <= 9'b101111000;
				8'b1101011: c <= 9'b11101111;
				8'b111100: c <= 9'b11011101;
				8'b1000111: c <= 9'b11011010;
				8'b1011111: c <= 9'b10001100;
				8'b1110100: c <= 9'b111;
				8'b101101: c <= 9'b10011001;
				8'b1010011: c <= 9'b100111;
				8'b1100001: c <= 9'b111011001;
				8'b110101: c <= 9'b1000111;
				8'b1000100: c <= 9'b101010101;
				8'b1010001: c <= 9'b100101110;
				8'b1010100: c <= 9'b110001110;
				8'b1100110: c <= 9'b101011001;
				8'b101010: c <= 9'b111110001;
				8'b1011110: c <= 9'b100;
				8'b1100111: c <= 9'b101111000;
				8'b1011010: c <= 9'b101111010;
				8'b1000010: c <= 9'b111001001;
				8'b111101: c <= 9'b11010;
				8'b110000: c <= 9'b1110011;
				8'b111110: c <= 9'b111100;
				8'b1100010: c <= 9'b110100111;
				8'b1110000: c <= 9'b100101011;
				8'b1101001: c <= 9'b11111101;
				8'b1110011: c <= 9'b11110101;
				8'b1001100: c <= 9'b10100110;
				8'b100001: c <= 9'b10010100;
				8'b1000110: c <= 9'b111101110;
				8'b1110010: c <= 9'b111101;
				8'b1010000: c <= 9'b101000101;
				8'b1111010: c <= 9'b101010101;
				8'b1010101: c <= 9'b101101100;
				8'b111011: c <= 9'b11111100;
				8'b1001101: c <= 9'b100101101;
				8'b111111: c <= 9'b1001110;
				8'b1101110: c <= 9'b100010110;
				8'b1111011: c <= 9'b10011100;
				8'b1001011: c <= 9'b110110011;
				8'b1101111: c <= 9'b110011000;
				8'b1101000: c <= 9'b1100000;
				8'b101100: c <= 9'b111000100;
				8'b100100: c <= 9'b111011001;
				8'b1111000: c <= 9'b10101010;
				8'b1000101: c <= 9'b101011110;
				8'b1011001: c <= 9'b11110010;
				8'b110100: c <= 9'b111011010;
				8'b1111001: c <= 9'b10001001;
				8'b1110001: c <= 9'b110001101;
				8'b1001111: c <= 9'b11100010;
				8'b1100101: c <= 9'b1011111;
				8'b1111110: c <= 9'b1010110;
				8'b1111100: c <= 9'b100001010;
				8'b1010110: c <= 9'b100000001;
				8'b110010: c <= 9'b1110010;
				8'b1101101: c <= 9'b100000111;
				8'b100011: c <= 9'b111111111;
				8'b1110101: c <= 9'b100001111;
				8'b1111101: c <= 9'b111011100;
				8'b101001: c <= 9'b111111101;
				8'b1010010: c <= 9'b10001100;
				8'b1011000: c <= 9'b1000000;
				8'b101110: c <= 9'b110000111;
				8'b1000001: c <= 9'b1000001;
				default: c <= 9'b0;
			endcase
			9'b1101011 : case(di)
				8'b1000011: c <= 9'b1110010;
				8'b101000: c <= 9'b101111000;
				8'b111010: c <= 9'b110101111;
				8'b110110: c <= 9'b111001110;
				8'b1100100: c <= 9'b1011100;
				8'b1000000: c <= 9'b110110011;
				8'b1110110: c <= 9'b11100100;
				8'b100101: c <= 9'b100001001;
				8'b101111: c <= 9'b1100011;
				8'b100110: c <= 9'b110001101;
				8'b1100011: c <= 9'b11101001;
				8'b1001000: c <= 9'b110111001;
				8'b111000: c <= 9'b110011110;
				8'b110001: c <= 9'b110110;
				8'b1010111: c <= 9'b100010;
				8'b1001110: c <= 9'b1100010;
				8'b1101010: c <= 9'b101101011;
				8'b1001001: c <= 9'b10011;
				8'b1100000: c <= 9'b101110100;
				8'b110111: c <= 9'b11011100;
				8'b1011101: c <= 9'b1101001;
				8'b1011011: c <= 9'b11101111;
				8'b111001: c <= 9'b110100010;
				8'b1001010: c <= 9'b101110011;
				8'b110011: c <= 9'b111010010;
				8'b1101100: c <= 9'b11110011;
				8'b1110111: c <= 9'b101000101;
				8'b101011: c <= 9'b111110101;
				8'b1101011: c <= 9'b10010101;
				8'b111100: c <= 9'b11011000;
				8'b1000111: c <= 9'b10110100;
				8'b1011111: c <= 9'b10111110;
				8'b1110100: c <= 9'b110101;
				8'b101101: c <= 9'b101110100;
				8'b1010011: c <= 9'b10000;
				8'b1100001: c <= 9'b10111001;
				8'b110101: c <= 9'b10001011;
				8'b1000100: c <= 9'b11000111;
				8'b1010001: c <= 9'b10;
				8'b1010100: c <= 9'b111101011;
				8'b1100110: c <= 9'b111001;
				8'b101010: c <= 9'b100100;
				8'b1011110: c <= 9'b100010;
				8'b1100111: c <= 9'b1011111;
				8'b1011010: c <= 9'b101100111;
				8'b1000010: c <= 9'b110111001;
				8'b111101: c <= 9'b100110110;
				8'b110000: c <= 9'b1000110;
				8'b111110: c <= 9'b11011;
				8'b1100010: c <= 9'b100010001;
				8'b1110000: c <= 9'b10;
				8'b1101001: c <= 9'b11110110;
				8'b1110011: c <= 9'b1111110;
				8'b1001100: c <= 9'b10001010;
				8'b100001: c <= 9'b100000111;
				8'b1000110: c <= 9'b11111;
				8'b1110010: c <= 9'b1000110;
				8'b1010000: c <= 9'b1100100;
				8'b1111010: c <= 9'b100000000;
				8'b1010101: c <= 9'b11011000;
				8'b111011: c <= 9'b101101111;
				8'b1001101: c <= 9'b110011111;
				8'b111111: c <= 9'b111111110;
				8'b1101110: c <= 9'b101111010;
				8'b1111011: c <= 9'b101010100;
				8'b1001011: c <= 9'b10010;
				8'b1101111: c <= 9'b11110;
				8'b1101000: c <= 9'b100100001;
				8'b101100: c <= 9'b11000000;
				8'b100100: c <= 9'b111110000;
				8'b1111000: c <= 9'b100111111;
				8'b1000101: c <= 9'b101100011;
				8'b1011001: c <= 9'b101010111;
				8'b110100: c <= 9'b111010000;
				8'b1111001: c <= 9'b1110100;
				8'b1110001: c <= 9'b11111010;
				8'b1001111: c <= 9'b101010110;
				8'b1100101: c <= 9'b111001110;
				8'b1111110: c <= 9'b1000100;
				8'b1111100: c <= 9'b110011110;
				8'b1010110: c <= 9'b101011011;
				8'b110010: c <= 9'b100111100;
				8'b1101101: c <= 9'b110110011;
				8'b100011: c <= 9'b100111;
				8'b1110101: c <= 9'b11110110;
				8'b1111101: c <= 9'b1011111;
				8'b101001: c <= 9'b100100000;
				8'b1010010: c <= 9'b101000101;
				8'b1011000: c <= 9'b1100110;
				8'b101110: c <= 9'b10010000;
				8'b1000001: c <= 9'b11000001;
				default: c <= 9'b0;
			endcase
			9'b111101011 : case(di)
				8'b1000011: c <= 9'b1010001;
				8'b101000: c <= 9'b100111;
				8'b111010: c <= 9'b100010;
				8'b110110: c <= 9'b110011011;
				8'b1100100: c <= 9'b1110101;
				8'b1000000: c <= 9'b1100000;
				8'b1110110: c <= 9'b100101010;
				8'b100101: c <= 9'b110110101;
				8'b101111: c <= 9'b1010011;
				8'b100110: c <= 9'b101011011;
				8'b1100011: c <= 9'b101001010;
				8'b1001000: c <= 9'b101000100;
				8'b111000: c <= 9'b101010111;
				8'b110001: c <= 9'b101001110;
				8'b1010111: c <= 9'b100010110;
				8'b1001110: c <= 9'b110010111;
				8'b1101010: c <= 9'b1011000;
				8'b1001001: c <= 9'b101101100;
				8'b1100000: c <= 9'b101001111;
				8'b110111: c <= 9'b10101111;
				8'b1011101: c <= 9'b110100011;
				8'b1011011: c <= 9'b111100;
				8'b111001: c <= 9'b1101111;
				8'b1001010: c <= 9'b10001000;
				8'b110011: c <= 9'b11111000;
				8'b1101100: c <= 9'b101110010;
				8'b1110111: c <= 9'b10100100;
				8'b101011: c <= 9'b101011;
				8'b1101011: c <= 9'b1011110;
				8'b111100: c <= 9'b111100;
				8'b1000111: c <= 9'b101001000;
				8'b1011111: c <= 9'b111111000;
				8'b1110100: c <= 9'b1000101;
				8'b101101: c <= 9'b1111111;
				8'b1010011: c <= 9'b10111101;
				8'b1100001: c <= 9'b10000110;
				8'b110101: c <= 9'b10101010;
				8'b1000100: c <= 9'b101011011;
				8'b1010001: c <= 9'b111011010;
				8'b1010100: c <= 9'b100011111;
				8'b1100110: c <= 9'b10100100;
				8'b101010: c <= 9'b1100010;
				8'b1011110: c <= 9'b100111;
				8'b1100111: c <= 9'b100011111;
				8'b1011010: c <= 9'b10101111;
				8'b1000010: c <= 9'b100100;
				8'b111101: c <= 9'b1011111;
				8'b110000: c <= 9'b101101000;
				8'b111110: c <= 9'b11100000;
				8'b1100010: c <= 9'b111101100;
				8'b1110000: c <= 9'b1001011;
				8'b1101001: c <= 9'b111110101;
				8'b1110011: c <= 9'b10100101;
				8'b1001100: c <= 9'b100110;
				8'b100001: c <= 9'b100011100;
				8'b1000110: c <= 9'b11101110;
				8'b1110010: c <= 9'b110000000;
				8'b1010000: c <= 9'b11010001;
				8'b1111010: c <= 9'b111111101;
				8'b1010101: c <= 9'b11011001;
				8'b111011: c <= 9'b110111010;
				8'b1001101: c <= 9'b10100100;
				8'b111111: c <= 9'b110000000;
				8'b1101110: c <= 9'b11001100;
				8'b1111011: c <= 9'b111;
				8'b1001011: c <= 9'b10000110;
				8'b1101111: c <= 9'b111010;
				8'b1101000: c <= 9'b10101101;
				8'b101100: c <= 9'b111101;
				8'b100100: c <= 9'b110010111;
				8'b1111000: c <= 9'b11101001;
				8'b1000101: c <= 9'b100100101;
				8'b1011001: c <= 9'b11110000;
				8'b110100: c <= 9'b111101100;
				8'b1111001: c <= 9'b100011;
				8'b1110001: c <= 9'b101110010;
				8'b1001111: c <= 9'b100100001;
				8'b1100101: c <= 9'b1000001;
				8'b1111110: c <= 9'b100111101;
				8'b1111100: c <= 9'b1111;
				8'b1010110: c <= 9'b111000010;
				8'b110010: c <= 9'b11010100;
				8'b1101101: c <= 9'b100011000;
				8'b100011: c <= 9'b101110100;
				8'b1110101: c <= 9'b101101001;
				8'b1111101: c <= 9'b1001100;
				8'b101001: c <= 9'b11000010;
				8'b1010010: c <= 9'b110100110;
				8'b1011000: c <= 9'b11110001;
				8'b101110: c <= 9'b101100011;
				8'b1000001: c <= 9'b101001;
				default: c <= 9'b0;
			endcase
			9'b11101110 : case(di)
				8'b1000011: c <= 9'b1100001;
				8'b101000: c <= 9'b111011101;
				8'b111010: c <= 9'b111100000;
				8'b110110: c <= 9'b11001001;
				8'b1100100: c <= 9'b101010100;
				8'b1000000: c <= 9'b101101110;
				8'b1110110: c <= 9'b101110110;
				8'b100101: c <= 9'b1001110;
				8'b101111: c <= 9'b10100110;
				8'b100110: c <= 9'b10110011;
				8'b1100011: c <= 9'b111011110;
				8'b1001000: c <= 9'b11111100;
				8'b111000: c <= 9'b110100000;
				8'b110001: c <= 9'b111111001;
				8'b1010111: c <= 9'b11000011;
				8'b1001110: c <= 9'b1111001;
				8'b1101010: c <= 9'b100100011;
				8'b1001001: c <= 9'b100000101;
				8'b1100000: c <= 9'b101111110;
				8'b110111: c <= 9'b110110000;
				8'b1011101: c <= 9'b100111000;
				8'b1011011: c <= 9'b111110001;
				8'b111001: c <= 9'b101111010;
				8'b1001010: c <= 9'b11100111;
				8'b110011: c <= 9'b1010000;
				8'b1101100: c <= 9'b111110011;
				8'b1110111: c <= 9'b10110011;
				8'b101011: c <= 9'b10101;
				8'b1101011: c <= 9'b101000100;
				8'b111100: c <= 9'b110000110;
				8'b1000111: c <= 9'b111111001;
				8'b1011111: c <= 9'b10100000;
				8'b1110100: c <= 9'b101111000;
				8'b101101: c <= 9'b1001000;
				8'b1010011: c <= 9'b11100;
				8'b1100001: c <= 9'b11000001;
				8'b110101: c <= 9'b10011111;
				8'b1000100: c <= 9'b100111000;
				8'b1010001: c <= 9'b111100010;
				8'b1010100: c <= 9'b1100111;
				8'b1100110: c <= 9'b111011011;
				8'b101010: c <= 9'b110100;
				8'b1011110: c <= 9'b100111101;
				8'b1100111: c <= 9'b11101101;
				8'b1011010: c <= 9'b111010100;
				8'b1000010: c <= 9'b110011110;
				8'b111101: c <= 9'b101100011;
				8'b110000: c <= 9'b10010110;
				8'b111110: c <= 9'b10001111;
				8'b1100010: c <= 9'b10011010;
				8'b1110000: c <= 9'b1100010;
				8'b1101001: c <= 9'b101110010;
				8'b1110011: c <= 9'b110101011;
				8'b1001100: c <= 9'b1111000;
				8'b100001: c <= 9'b11100011;
				8'b1000110: c <= 9'b10101001;
				8'b1110010: c <= 9'b1100100;
				8'b1010000: c <= 9'b111101000;
				8'b1111010: c <= 9'b101110100;
				8'b1010101: c <= 9'b111100101;
				8'b111011: c <= 9'b110010101;
				8'b1001101: c <= 9'b110010111;
				8'b111111: c <= 9'b11110000;
				8'b1101110: c <= 9'b11000001;
				8'b1111011: c <= 9'b101111011;
				8'b1001011: c <= 9'b111011110;
				8'b1101111: c <= 9'b10100100;
				8'b1101000: c <= 9'b111111010;
				8'b101100: c <= 9'b10100;
				8'b100100: c <= 9'b101111000;
				8'b1111000: c <= 9'b100100011;
				8'b1000101: c <= 9'b1110001;
				8'b1011001: c <= 9'b101001000;
				8'b110100: c <= 9'b10000000;
				8'b1111001: c <= 9'b1101101;
				8'b1110001: c <= 9'b11000111;
				8'b1001111: c <= 9'b111100100;
				8'b1100101: c <= 9'b100110101;
				8'b1111110: c <= 9'b11100101;
				8'b1111100: c <= 9'b10000110;
				8'b1010110: c <= 9'b110100101;
				8'b110010: c <= 9'b111011101;
				8'b1101101: c <= 9'b101001011;
				8'b100011: c <= 9'b111111;
				8'b1110101: c <= 9'b10011010;
				8'b1111101: c <= 9'b100110000;
				8'b101001: c <= 9'b11001;
				8'b1010010: c <= 9'b110010110;
				8'b1011000: c <= 9'b11011011;
				8'b101110: c <= 9'b101001111;
				8'b1000001: c <= 9'b101011101;
				default: c <= 9'b0;
			endcase
			9'b101111011 : case(di)
				8'b1000011: c <= 9'b111011110;
				8'b101000: c <= 9'b11001010;
				8'b111010: c <= 9'b101000111;
				8'b110110: c <= 9'b11100011;
				8'b1100100: c <= 9'b101110010;
				8'b1000000: c <= 9'b100010010;
				8'b1110110: c <= 9'b10000;
				8'b100101: c <= 9'b10100110;
				8'b101111: c <= 9'b11101;
				8'b100110: c <= 9'b11110000;
				8'b1100011: c <= 9'b110100101;
				8'b1001000: c <= 9'b11000000;
				8'b111000: c <= 9'b10011011;
				8'b110001: c <= 9'b11001001;
				8'b1010111: c <= 9'b1001111;
				8'b1001110: c <= 9'b110001001;
				8'b1101010: c <= 9'b111011011;
				8'b1001001: c <= 9'b111110;
				8'b1100000: c <= 9'b100000101;
				8'b110111: c <= 9'b111000011;
				8'b1011101: c <= 9'b111101000;
				8'b1011011: c <= 9'b1000100;
				8'b111001: c <= 9'b111111101;
				8'b1001010: c <= 9'b111101101;
				8'b110011: c <= 9'b11110010;
				8'b1101100: c <= 9'b1111000;
				8'b1110111: c <= 9'b100000011;
				8'b101011: c <= 9'b100010001;
				8'b1101011: c <= 9'b111110000;
				8'b111100: c <= 9'b11101100;
				8'b1000111: c <= 9'b1111001;
				8'b1011111: c <= 9'b111101010;
				8'b1110100: c <= 9'b101101111;
				8'b101101: c <= 9'b101101000;
				8'b1010011: c <= 9'b100100101;
				8'b1100001: c <= 9'b111100110;
				8'b110101: c <= 9'b110111;
				8'b1000100: c <= 9'b111101111;
				8'b1010001: c <= 9'b111010100;
				8'b1010100: c <= 9'b1111101;
				8'b1100110: c <= 9'b10101101;
				8'b101010: c <= 9'b110101001;
				8'b1011110: c <= 9'b11100000;
				8'b1100111: c <= 9'b1101110;
				8'b1011010: c <= 9'b1110011;
				8'b1000010: c <= 9'b1000010;
				8'b111101: c <= 9'b1100101;
				8'b110000: c <= 9'b11011;
				8'b111110: c <= 9'b111000110;
				8'b1100010: c <= 9'b10100000;
				8'b1110000: c <= 9'b11101001;
				8'b1101001: c <= 9'b111010111;
				8'b1110011: c <= 9'b11010;
				8'b1001100: c <= 9'b10110011;
				8'b100001: c <= 9'b1100101;
				8'b1000110: c <= 9'b10010101;
				8'b1110010: c <= 9'b101011001;
				8'b1010000: c <= 9'b11100001;
				8'b1111010: c <= 9'b100000101;
				8'b1010101: c <= 9'b111101100;
				8'b111011: c <= 9'b100001010;
				8'b1001101: c <= 9'b111001010;
				8'b111111: c <= 9'b100011001;
				8'b1101110: c <= 9'b1111;
				8'b1111011: c <= 9'b1111;
				8'b1001011: c <= 9'b101010111;
				8'b1101111: c <= 9'b110111110;
				8'b1101000: c <= 9'b11010011;
				8'b101100: c <= 9'b100110100;
				8'b100100: c <= 9'b1100100;
				8'b1111000: c <= 9'b100101;
				8'b1000101: c <= 9'b10100000;
				8'b1011001: c <= 9'b1;
				8'b110100: c <= 9'b101010110;
				8'b1111001: c <= 9'b11101111;
				8'b1110001: c <= 9'b11000;
				8'b1001111: c <= 9'b10101111;
				8'b1100101: c <= 9'b111000;
				8'b1111110: c <= 9'b100101110;
				8'b1111100: c <= 9'b110001000;
				8'b1010110: c <= 9'b10001111;
				8'b110010: c <= 9'b101000110;
				8'b1101101: c <= 9'b10111010;
				8'b100011: c <= 9'b10000110;
				8'b1110101: c <= 9'b11100100;
				8'b1111101: c <= 9'b10010001;
				8'b101001: c <= 9'b111101010;
				8'b1010010: c <= 9'b10101011;
				8'b1011000: c <= 9'b11010011;
				8'b101110: c <= 9'b110110110;
				8'b1000001: c <= 9'b101000110;
				default: c <= 9'b0;
			endcase
			9'b111110 : case(di)
				8'b1000011: c <= 9'b101100111;
				8'b101000: c <= 9'b110101101;
				8'b111010: c <= 9'b10110110;
				8'b110110: c <= 9'b11011110;
				8'b1100100: c <= 9'b10101100;
				8'b1000000: c <= 9'b100000000;
				8'b1110110: c <= 9'b111110110;
				8'b100101: c <= 9'b1110;
				8'b101111: c <= 9'b11001100;
				8'b100110: c <= 9'b10100101;
				8'b1100011: c <= 9'b11111100;
				8'b1001000: c <= 9'b10100011;
				8'b111000: c <= 9'b100011111;
				8'b110001: c <= 9'b11000010;
				8'b1010111: c <= 9'b1000100;
				8'b1001110: c <= 9'b11100000;
				8'b1101010: c <= 9'b110110101;
				8'b1001001: c <= 9'b101010010;
				8'b1100000: c <= 9'b100111000;
				8'b110111: c <= 9'b110100100;
				8'b1011101: c <= 9'b101111000;
				8'b1011011: c <= 9'b110101101;
				8'b111001: c <= 9'b101001011;
				8'b1001010: c <= 9'b101000010;
				8'b110011: c <= 9'b1110111;
				8'b1101100: c <= 9'b101100100;
				8'b1110111: c <= 9'b110101110;
				8'b101011: c <= 9'b11100000;
				8'b1101011: c <= 9'b111010000;
				8'b111100: c <= 9'b100101;
				8'b1000111: c <= 9'b101110101;
				8'b1011111: c <= 9'b10011110;
				8'b1110100: c <= 9'b10101100;
				8'b101101: c <= 9'b101010;
				8'b1010011: c <= 9'b10011010;
				8'b1100001: c <= 9'b11001110;
				8'b110101: c <= 9'b11011100;
				8'b1000100: c <= 9'b111001110;
				8'b1010001: c <= 9'b1001010;
				8'b1010100: c <= 9'b111111110;
				8'b1100110: c <= 9'b10101101;
				8'b101010: c <= 9'b110100010;
				8'b1011110: c <= 9'b111010000;
				8'b1100111: c <= 9'b100100000;
				8'b1011010: c <= 9'b110110111;
				8'b1000010: c <= 9'b100100010;
				8'b111101: c <= 9'b10010;
				8'b110000: c <= 9'b11110110;
				8'b111110: c <= 9'b111011010;
				8'b1100010: c <= 9'b1001011;
				8'b1110000: c <= 9'b100011101;
				8'b1101001: c <= 9'b1010000;
				8'b1110011: c <= 9'b1010001;
				8'b1001100: c <= 9'b11011110;
				8'b100001: c <= 9'b1010001;
				8'b1000110: c <= 9'b111001010;
				8'b1110010: c <= 9'b1011110;
				8'b1010000: c <= 9'b11011000;
				8'b1111010: c <= 9'b11100000;
				8'b1010101: c <= 9'b11011010;
				8'b111011: c <= 9'b101100001;
				8'b1001101: c <= 9'b100101100;
				8'b111111: c <= 9'b111010010;
				8'b1101110: c <= 9'b110000;
				8'b1111011: c <= 9'b110110101;
				8'b1001011: c <= 9'b101001100;
				8'b1101111: c <= 9'b101010111;
				8'b1101000: c <= 9'b110011010;
				8'b101100: c <= 9'b101100110;
				8'b100100: c <= 9'b110100111;
				8'b1111000: c <= 9'b10111001;
				8'b1000101: c <= 9'b10001000;
				8'b1011001: c <= 9'b110100101;
				8'b110100: c <= 9'b1110011;
				8'b1111001: c <= 9'b1111001;
				8'b1110001: c <= 9'b10110110;
				8'b1001111: c <= 9'b11000;
				8'b1100101: c <= 9'b110111;
				8'b1111110: c <= 9'b110110100;
				8'b1111100: c <= 9'b111010;
				8'b1010110: c <= 9'b111000111;
				8'b110010: c <= 9'b1011110;
				8'b1101101: c <= 9'b110111100;
				8'b100011: c <= 9'b1000011;
				8'b1110101: c <= 9'b100010011;
				8'b1111101: c <= 9'b110100101;
				8'b101001: c <= 9'b10000110;
				8'b1010010: c <= 9'b111011010;
				8'b1011000: c <= 9'b11111100;
				8'b101110: c <= 9'b10100110;
				8'b1000001: c <= 9'b100111;
				default: c <= 9'b0;
			endcase
			9'b10011110 : case(di)
				8'b1000011: c <= 9'b1101100;
				8'b101000: c <= 9'b101100000;
				8'b111010: c <= 9'b100011000;
				8'b110110: c <= 9'b111101010;
				8'b1100100: c <= 9'b110001100;
				8'b1000000: c <= 9'b101110000;
				8'b1110110: c <= 9'b111000011;
				8'b100101: c <= 9'b110101010;
				8'b101111: c <= 9'b10111100;
				8'b100110: c <= 9'b110111100;
				8'b1100011: c <= 9'b100011000;
				8'b1001000: c <= 9'b110001010;
				8'b111000: c <= 9'b11001101;
				8'b110001: c <= 9'b111010010;
				8'b1010111: c <= 9'b111101101;
				8'b1001110: c <= 9'b100010111;
				8'b1101010: c <= 9'b1000011;
				8'b1001001: c <= 9'b101111000;
				8'b1100000: c <= 9'b1100101;
				8'b110111: c <= 9'b111000;
				8'b1011101: c <= 9'b11100110;
				8'b1011011: c <= 9'b10010111;
				8'b111001: c <= 9'b100110010;
				8'b1001010: c <= 9'b100111111;
				8'b110011: c <= 9'b10011010;
				8'b1101100: c <= 9'b111011010;
				8'b1110111: c <= 9'b111100;
				8'b101011: c <= 9'b100110010;
				8'b1101011: c <= 9'b101011011;
				8'b111100: c <= 9'b110110011;
				8'b1000111: c <= 9'b10001011;
				8'b1011111: c <= 9'b10100011;
				8'b1110100: c <= 9'b110100001;
				8'b101101: c <= 9'b110001010;
				8'b1010011: c <= 9'b10110111;
				8'b1100001: c <= 9'b10110010;
				8'b110101: c <= 9'b111101001;
				8'b1000100: c <= 9'b100011100;
				8'b1010001: c <= 9'b111100000;
				8'b1010100: c <= 9'b100101101;
				8'b1100110: c <= 9'b11000000;
				8'b101010: c <= 9'b100001101;
				8'b1011110: c <= 9'b111001100;
				8'b1100111: c <= 9'b100010101;
				8'b1011010: c <= 9'b1101111;
				8'b1000010: c <= 9'b101010001;
				8'b111101: c <= 9'b100110101;
				8'b110000: c <= 9'b1010011;
				8'b111110: c <= 9'b10000101;
				8'b1100010: c <= 9'b10;
				8'b1110000: c <= 9'b10000011;
				8'b1101001: c <= 9'b111001000;
				8'b1110011: c <= 9'b100010110;
				8'b1001100: c <= 9'b101100011;
				8'b100001: c <= 9'b110010010;
				8'b1000110: c <= 9'b11100110;
				8'b1110010: c <= 9'b101011;
				8'b1010000: c <= 9'b111101100;
				8'b1111010: c <= 9'b100011000;
				8'b1010101: c <= 9'b100001110;
				8'b111011: c <= 9'b100000010;
				8'b1001101: c <= 9'b10001100;
				8'b111111: c <= 9'b111011111;
				8'b1101110: c <= 9'b11110;
				8'b1111011: c <= 9'b110010001;
				8'b1001011: c <= 9'b11000;
				8'b1101111: c <= 9'b101110001;
				8'b1101000: c <= 9'b111000001;
				8'b101100: c <= 9'b111101101;
				8'b100100: c <= 9'b101100111;
				8'b1111000: c <= 9'b100010000;
				8'b1000101: c <= 9'b11100001;
				8'b1011001: c <= 9'b11111101;
				8'b110100: c <= 9'b1111000;
				8'b1111001: c <= 9'b100100101;
				8'b1110001: c <= 9'b110111;
				8'b1001111: c <= 9'b110011010;
				8'b1100101: c <= 9'b101111000;
				8'b1111110: c <= 9'b11110101;
				8'b1111100: c <= 9'b100011001;
				8'b1010110: c <= 9'b10101101;
				8'b110010: c <= 9'b101100;
				8'b1101101: c <= 9'b101001100;
				8'b100011: c <= 9'b10101011;
				8'b1110101: c <= 9'b111100101;
				8'b1111101: c <= 9'b110110111;
				8'b101001: c <= 9'b11000001;
				8'b1010010: c <= 9'b10011001;
				8'b1011000: c <= 9'b1011111;
				8'b101110: c <= 9'b110110111;
				8'b1000001: c <= 9'b111011011;
				default: c <= 9'b0;
			endcase
			9'b111000001 : case(di)
				8'b1000011: c <= 9'b10111111;
				8'b101000: c <= 9'b111011101;
				8'b111010: c <= 9'b11010001;
				8'b110110: c <= 9'b111100011;
				8'b1100100: c <= 9'b11100001;
				8'b1000000: c <= 9'b1010001;
				8'b1110110: c <= 9'b1100100;
				8'b100101: c <= 9'b11111100;
				8'b101111: c <= 9'b110011011;
				8'b100110: c <= 9'b101110101;
				8'b1100011: c <= 9'b110111001;
				8'b1001000: c <= 9'b100101101;
				8'b111000: c <= 9'b11100001;
				8'b110001: c <= 9'b111100011;
				8'b1010111: c <= 9'b1100000;
				8'b1001110: c <= 9'b1011;
				8'b1101010: c <= 9'b11111101;
				8'b1001001: c <= 9'b111100001;
				8'b1100000: c <= 9'b100000101;
				8'b110111: c <= 9'b110001111;
				8'b1011101: c <= 9'b110100110;
				8'b1011011: c <= 9'b100100111;
				8'b111001: c <= 9'b100011100;
				8'b1001010: c <= 9'b110110010;
				8'b110011: c <= 9'b1100000;
				8'b1101100: c <= 9'b100100110;
				8'b1110111: c <= 9'b11001101;
				8'b101011: c <= 9'b110110100;
				8'b1101011: c <= 9'b10110100;
				8'b111100: c <= 9'b110011111;
				8'b1000111: c <= 9'b11001100;
				8'b1011111: c <= 9'b1011100;
				8'b1110100: c <= 9'b1111011;
				8'b101101: c <= 9'b100100011;
				8'b1010011: c <= 9'b10111101;
				8'b1100001: c <= 9'b101010;
				8'b110101: c <= 9'b10111010;
				8'b1000100: c <= 9'b1000011;
				8'b1010001: c <= 9'b1101;
				8'b1010100: c <= 9'b1110010;
				8'b1100110: c <= 9'b11110100;
				8'b101010: c <= 9'b100100;
				8'b1011110: c <= 9'b10101011;
				8'b1100111: c <= 9'b110111111;
				8'b1011010: c <= 9'b11010111;
				8'b1000010: c <= 9'b110100000;
				8'b111101: c <= 9'b11100100;
				8'b110000: c <= 9'b11010110;
				8'b111110: c <= 9'b111;
				8'b1100010: c <= 9'b100100001;
				8'b1110000: c <= 9'b110100110;
				8'b1101001: c <= 9'b10000000;
				8'b1110011: c <= 9'b10001100;
				8'b1001100: c <= 9'b1010011;
				8'b100001: c <= 9'b10010011;
				8'b1000110: c <= 9'b100101010;
				8'b1110010: c <= 9'b100000001;
				8'b1010000: c <= 9'b11000110;
				8'b1111010: c <= 9'b101100010;
				8'b1010101: c <= 9'b111110101;
				8'b111011: c <= 9'b10011001;
				8'b1001101: c <= 9'b111010111;
				8'b111111: c <= 9'b10011;
				8'b1101110: c <= 9'b101011010;
				8'b1111011: c <= 9'b11010111;
				8'b1001011: c <= 9'b10001000;
				8'b1101111: c <= 9'b11011;
				8'b1101000: c <= 9'b10110110;
				8'b101100: c <= 9'b1101;
				8'b100100: c <= 9'b101100100;
				8'b1111000: c <= 9'b101101001;
				8'b1000101: c <= 9'b11010100;
				8'b1011001: c <= 9'b111111101;
				8'b110100: c <= 9'b100111100;
				8'b1111001: c <= 9'b10101111;
				8'b1110001: c <= 9'b111010;
				8'b1001111: c <= 9'b110100101;
				8'b1100101: c <= 9'b101101110;
				8'b1111110: c <= 9'b11011001;
				8'b1111100: c <= 9'b111001;
				8'b1010110: c <= 9'b111111111;
				8'b110010: c <= 9'b100101111;
				8'b1101101: c <= 9'b111111000;
				8'b100011: c <= 9'b111001010;
				8'b1110101: c <= 9'b1110111;
				8'b1111101: c <= 9'b101111110;
				8'b101001: c <= 9'b10011100;
				8'b1010010: c <= 9'b1110010;
				8'b1011000: c <= 9'b101101011;
				8'b101110: c <= 9'b10100011;
				8'b1000001: c <= 9'b100010010;
				default: c <= 9'b0;
			endcase
			9'b11010110 : case(di)
				8'b1000011: c <= 9'b111011011;
				8'b101000: c <= 9'b110001;
				8'b111010: c <= 9'b1111101;
				8'b110110: c <= 9'b110000111;
				8'b1100100: c <= 9'b100101000;
				8'b1000000: c <= 9'b111110001;
				8'b1110110: c <= 9'b11010010;
				8'b100101: c <= 9'b10001110;
				8'b101111: c <= 9'b10100;
				8'b100110: c <= 9'b100000011;
				8'b1100011: c <= 9'b11001000;
				8'b1001000: c <= 9'b11011100;
				8'b111000: c <= 9'b10010101;
				8'b110001: c <= 9'b100001001;
				8'b1010111: c <= 9'b10010011;
				8'b1001110: c <= 9'b111000011;
				8'b1101010: c <= 9'b10110011;
				8'b1001001: c <= 9'b110110110;
				8'b1100000: c <= 9'b101101100;
				8'b110111: c <= 9'b111001010;
				8'b1011101: c <= 9'b110111000;
				8'b1011011: c <= 9'b1011100;
				8'b111001: c <= 9'b10110011;
				8'b1001010: c <= 9'b1101000;
				8'b110011: c <= 9'b100001111;
				8'b1101100: c <= 9'b10011001;
				8'b1110111: c <= 9'b101101100;
				8'b101011: c <= 9'b100011011;
				8'b1101011: c <= 9'b10;
				8'b111100: c <= 9'b1000110;
				8'b1000111: c <= 9'b100010000;
				8'b1011111: c <= 9'b101010001;
				8'b1110100: c <= 9'b100111101;
				8'b101101: c <= 9'b101001111;
				8'b1010011: c <= 9'b110000010;
				8'b1100001: c <= 9'b110110010;
				8'b110101: c <= 9'b1111111;
				8'b1000100: c <= 9'b1000001;
				8'b1010001: c <= 9'b11010100;
				8'b1010100: c <= 9'b1110101;
				8'b1100110: c <= 9'b101100010;
				8'b101010: c <= 9'b1010000;
				8'b1011110: c <= 9'b101110000;
				8'b1100111: c <= 9'b110101010;
				8'b1011010: c <= 9'b111001110;
				8'b1000010: c <= 9'b101;
				8'b111101: c <= 9'b10001101;
				8'b110000: c <= 9'b1100100;
				8'b111110: c <= 9'b11;
				8'b1100010: c <= 9'b11111011;
				8'b1110000: c <= 9'b10000100;
				8'b1101001: c <= 9'b110010;
				8'b1110011: c <= 9'b11010111;
				8'b1001100: c <= 9'b100010000;
				8'b100001: c <= 9'b1000000;
				8'b1000110: c <= 9'b11100110;
				8'b1110010: c <= 9'b10100110;
				8'b1010000: c <= 9'b111001000;
				8'b1111010: c <= 9'b100111110;
				8'b1010101: c <= 9'b100111110;
				8'b111011: c <= 9'b111110000;
				8'b1001101: c <= 9'b10110111;
				8'b111111: c <= 9'b100011111;
				8'b1101110: c <= 9'b10110111;
				8'b1111011: c <= 9'b1101100;
				8'b1001011: c <= 9'b100101101;
				8'b1101111: c <= 9'b11001;
				8'b1101000: c <= 9'b110101111;
				8'b101100: c <= 9'b1111000;
				8'b100100: c <= 9'b11001000;
				8'b1111000: c <= 9'b11111011;
				8'b1000101: c <= 9'b1011010;
				8'b1011001: c <= 9'b100100111;
				8'b110100: c <= 9'b110010101;
				8'b1111001: c <= 9'b11010101;
				8'b1110001: c <= 9'b110011111;
				8'b1001111: c <= 9'b111000;
				8'b1100101: c <= 9'b110110;
				8'b1111110: c <= 9'b10010011;
				8'b1111100: c <= 9'b111101111;
				8'b1010110: c <= 9'b11000011;
				8'b110010: c <= 9'b101100100;
				8'b1101101: c <= 9'b1001010;
				8'b100011: c <= 9'b111001011;
				8'b1110101: c <= 9'b11110;
				8'b1111101: c <= 9'b11000100;
				8'b101001: c <= 9'b10100110;
				8'b1010010: c <= 9'b10000111;
				8'b1011000: c <= 9'b110001111;
				8'b101110: c <= 9'b110110100;
				8'b1000001: c <= 9'b101101101;
				default: c <= 9'b0;
			endcase
			9'b10000100 : case(di)
				8'b1000011: c <= 9'b101011110;
				8'b101000: c <= 9'b110010010;
				8'b111010: c <= 9'b101100000;
				8'b110110: c <= 9'b11111010;
				8'b1100100: c <= 9'b1000011;
				8'b1000000: c <= 9'b100000001;
				8'b1110110: c <= 9'b101110001;
				8'b100101: c <= 9'b110110010;
				8'b101111: c <= 9'b10110;
				8'b100110: c <= 9'b100010101;
				8'b1100011: c <= 9'b101100001;
				8'b1001000: c <= 9'b110100101;
				8'b111000: c <= 9'b11000001;
				8'b110001: c <= 9'b1001;
				8'b1010111: c <= 9'b110110110;
				8'b1001110: c <= 9'b10001010;
				8'b1101010: c <= 9'b10011000;
				8'b1001001: c <= 9'b111111110;
				8'b1100000: c <= 9'b10101101;
				8'b110111: c <= 9'b100011010;
				8'b1011101: c <= 9'b11100100;
				8'b1011011: c <= 9'b1111010;
				8'b111001: c <= 9'b10100011;
				8'b1001010: c <= 9'b100110110;
				8'b110011: c <= 9'b100011110;
				8'b1101100: c <= 9'b100000010;
				8'b1110111: c <= 9'b110010001;
				8'b101011: c <= 9'b111101000;
				8'b1101011: c <= 9'b110110011;
				8'b111100: c <= 9'b101001000;
				8'b1000111: c <= 9'b11101;
				8'b1011111: c <= 9'b10011;
				8'b1110100: c <= 9'b10111000;
				8'b101101: c <= 9'b100111011;
				8'b1010011: c <= 9'b10001000;
				8'b1100001: c <= 9'b110010110;
				8'b110101: c <= 9'b1011011;
				8'b1000100: c <= 9'b101010;
				8'b1010001: c <= 9'b11001101;
				8'b1010100: c <= 9'b10111110;
				8'b1100110: c <= 9'b101101100;
				8'b101010: c <= 9'b111000011;
				8'b1011110: c <= 9'b10110110;
				8'b1100111: c <= 9'b111000111;
				8'b1011010: c <= 9'b111100010;
				8'b1000010: c <= 9'b110100;
				8'b111101: c <= 9'b11011100;
				8'b110000: c <= 9'b101110101;
				8'b111110: c <= 9'b111011001;
				8'b1100010: c <= 9'b100111;
				8'b1110000: c <= 9'b100000011;
				8'b1101001: c <= 9'b11001101;
				8'b1110011: c <= 9'b10011001;
				8'b1001100: c <= 9'b101101001;
				8'b100001: c <= 9'b110000110;
				8'b1000110: c <= 9'b110011010;
				8'b1110010: c <= 9'b1101010;
				8'b1010000: c <= 9'b11001;
				8'b1111010: c <= 9'b1111011;
				8'b1010101: c <= 9'b101100;
				8'b111011: c <= 9'b101100100;
				8'b1001101: c <= 9'b111100000;
				8'b111111: c <= 9'b10110111;
				8'b1101110: c <= 9'b111011010;
				8'b1111011: c <= 9'b11110111;
				8'b1001011: c <= 9'b10010101;
				8'b1101111: c <= 9'b10001000;
				8'b1101000: c <= 9'b110011010;
				8'b101100: c <= 9'b11100000;
				8'b100100: c <= 9'b1011;
				8'b1111000: c <= 9'b10001100;
				8'b1000101: c <= 9'b10011011;
				8'b1011001: c <= 9'b101011000;
				8'b110100: c <= 9'b101101101;
				8'b1111001: c <= 9'b101110;
				8'b1110001: c <= 9'b1101000;
				8'b1001111: c <= 9'b100000101;
				8'b1100101: c <= 9'b1011;
				8'b1111110: c <= 9'b1101;
				8'b1111100: c <= 9'b111010110;
				8'b1010110: c <= 9'b1110101;
				8'b110010: c <= 9'b101011;
				8'b1101101: c <= 9'b1001000;
				8'b100011: c <= 9'b101110101;
				8'b1110101: c <= 9'b101101100;
				8'b1111101: c <= 9'b11000100;
				8'b101001: c <= 9'b10100101;
				8'b1010010: c <= 9'b11110000;
				8'b1011000: c <= 9'b100010111;
				8'b101110: c <= 9'b101100;
				8'b1000001: c <= 9'b10011;
				default: c <= 9'b0;
			endcase
			9'b100011110 : case(di)
				8'b1000011: c <= 9'b100110;
				8'b101000: c <= 9'b101100101;
				8'b111010: c <= 9'b10111000;
				8'b110110: c <= 9'b11000111;
				8'b1100100: c <= 9'b11001011;
				8'b1000000: c <= 9'b11010101;
				8'b1110110: c <= 9'b1011100;
				8'b100101: c <= 9'b11100010;
				8'b101111: c <= 9'b100101111;
				8'b100110: c <= 9'b1011111;
				8'b1100011: c <= 9'b1101010;
				8'b1001000: c <= 9'b101101001;
				8'b111000: c <= 9'b111100000;
				8'b110001: c <= 9'b100011101;
				8'b1010111: c <= 9'b100101001;
				8'b1001110: c <= 9'b111010010;
				8'b1101010: c <= 9'b1111111;
				8'b1001001: c <= 9'b101011110;
				8'b1100000: c <= 9'b110;
				8'b110111: c <= 9'b110001101;
				8'b1011101: c <= 9'b100100111;
				8'b1011011: c <= 9'b111100101;
				8'b111001: c <= 9'b11010111;
				8'b1001010: c <= 9'b10101011;
				8'b110011: c <= 9'b100011000;
				8'b1101100: c <= 9'b10001111;
				8'b1110111: c <= 9'b110110110;
				8'b101011: c <= 9'b1000011;
				8'b1101011: c <= 9'b11100101;
				8'b111100: c <= 9'b111011010;
				8'b1000111: c <= 9'b110110;
				8'b1011111: c <= 9'b100110001;
				8'b1110100: c <= 9'b110011100;
				8'b101101: c <= 9'b100000100;
				8'b1010011: c <= 9'b1110011;
				8'b1100001: c <= 9'b110000101;
				8'b110101: c <= 9'b100000111;
				8'b1000100: c <= 9'b110110000;
				8'b1010001: c <= 9'b1001010;
				8'b1010100: c <= 9'b11100;
				8'b1100110: c <= 9'b111000101;
				8'b101010: c <= 9'b100111010;
				8'b1011110: c <= 9'b111010000;
				8'b1100111: c <= 9'b10001001;
				8'b1011010: c <= 9'b11111000;
				8'b1000010: c <= 9'b101111010;
				8'b111101: c <= 9'b110101011;
				8'b110000: c <= 9'b110011100;
				8'b111110: c <= 9'b10110100;
				8'b1100010: c <= 9'b110010100;
				8'b1110000: c <= 9'b111001101;
				8'b1101001: c <= 9'b100101111;
				8'b1110011: c <= 9'b101100110;
				8'b1001100: c <= 9'b101001110;
				8'b100001: c <= 9'b100001101;
				8'b1000110: c <= 9'b11110110;
				8'b1110010: c <= 9'b101001111;
				8'b1010000: c <= 9'b11101101;
				8'b1111010: c <= 9'b10111;
				8'b1010101: c <= 9'b111001101;
				8'b111011: c <= 9'b110010010;
				8'b1001101: c <= 9'b11110;
				8'b111111: c <= 9'b100011001;
				8'b1101110: c <= 9'b110011011;
				8'b1111011: c <= 9'b11110111;
				8'b1001011: c <= 9'b11011011;
				8'b1101111: c <= 9'b10010011;
				8'b1101000: c <= 9'b110001111;
				8'b101100: c <= 9'b1101100;
				8'b100100: c <= 9'b11010010;
				8'b1111000: c <= 9'b111000111;
				8'b1000101: c <= 9'b10010011;
				8'b1011001: c <= 9'b1100;
				8'b110100: c <= 9'b1111;
				8'b1111001: c <= 9'b1000101;
				8'b1110001: c <= 9'b1000010;
				8'b1001111: c <= 9'b1100111;
				8'b1100101: c <= 9'b100010001;
				8'b1111110: c <= 9'b101011010;
				8'b1111100: c <= 9'b10010;
				8'b1010110: c <= 9'b110000111;
				8'b110010: c <= 9'b110011;
				8'b1101101: c <= 9'b11111011;
				8'b100011: c <= 9'b11000111;
				8'b1110101: c <= 9'b100010111;
				8'b1111101: c <= 9'b100111100;
				8'b101001: c <= 9'b101011;
				8'b1010010: c <= 9'b10110101;
				8'b1011000: c <= 9'b1001001;
				8'b101110: c <= 9'b100011100;
				8'b1000001: c <= 9'b111;
				default: c <= 9'b0;
			endcase
			9'b100110001 : case(di)
				8'b1000011: c <= 9'b101100;
				8'b101000: c <= 9'b1101111;
				8'b111010: c <= 9'b11000010;
				8'b110110: c <= 9'b11111010;
				8'b1100100: c <= 9'b10101000;
				8'b1000000: c <= 9'b10111000;
				8'b1110110: c <= 9'b10010011;
				8'b100101: c <= 9'b11001010;
				8'b101111: c <= 9'b100110110;
				8'b100110: c <= 9'b11110010;
				8'b1100011: c <= 9'b10011111;
				8'b1001000: c <= 9'b10001110;
				8'b111000: c <= 9'b100111110;
				8'b110001: c <= 9'b1;
				8'b1010111: c <= 9'b10110001;
				8'b1001110: c <= 9'b10111110;
				8'b1101010: c <= 9'b101000010;
				8'b1001001: c <= 9'b100011100;
				8'b1100000: c <= 9'b101101000;
				8'b110111: c <= 9'b110100011;
				8'b1011101: c <= 9'b10100011;
				8'b1011011: c <= 9'b111101000;
				8'b111001: c <= 9'b110010111;
				8'b1001010: c <= 9'b11001010;
				8'b110011: c <= 9'b111;
				8'b1101100: c <= 9'b111001011;
				8'b1110111: c <= 9'b101000001;
				8'b101011: c <= 9'b10101001;
				8'b1101011: c <= 9'b110010100;
				8'b111100: c <= 9'b101010001;
				8'b1000111: c <= 9'b10001010;
				8'b1011111: c <= 9'b110010;
				8'b1110100: c <= 9'b101110000;
				8'b101101: c <= 9'b100000011;
				8'b1010011: c <= 9'b11101000;
				8'b1100001: c <= 9'b10101111;
				8'b110101: c <= 9'b110011001;
				8'b1000100: c <= 9'b110011001;
				8'b1010001: c <= 9'b10011101;
				8'b1010100: c <= 9'b10101111;
				8'b1100110: c <= 9'b1101100;
				8'b101010: c <= 9'b11100001;
				8'b1011110: c <= 9'b1001001;
				8'b1100111: c <= 9'b110001110;
				8'b1011010: c <= 9'b100011010;
				8'b1000010: c <= 9'b111001001;
				8'b111101: c <= 9'b101100011;
				8'b110000: c <= 9'b11010010;
				8'b111110: c <= 9'b10100010;
				8'b1100010: c <= 9'b110100010;
				8'b1110000: c <= 9'b1001000;
				8'b1101001: c <= 9'b10101000;
				8'b1110011: c <= 9'b110011;
				8'b1001100: c <= 9'b10111;
				8'b100001: c <= 9'b100110110;
				8'b1000110: c <= 9'b10001111;
				8'b1110010: c <= 9'b111010010;
				8'b1010000: c <= 9'b101110100;
				8'b1111010: c <= 9'b101001;
				8'b1010101: c <= 9'b10000011;
				8'b111011: c <= 9'b100101;
				8'b1001101: c <= 9'b1100100;
				8'b111111: c <= 9'b110100010;
				8'b1101110: c <= 9'b11101001;
				8'b1111011: c <= 9'b101110110;
				8'b1001011: c <= 9'b100111100;
				8'b1101111: c <= 9'b110001100;
				8'b1101000: c <= 9'b10011011;
				8'b101100: c <= 9'b110100111;
				8'b100100: c <= 9'b11011;
				8'b1111000: c <= 9'b11100010;
				8'b1000101: c <= 9'b111001010;
				8'b1011001: c <= 9'b1101001;
				8'b110100: c <= 9'b1001001;
				8'b1111001: c <= 9'b101111100;
				8'b1110001: c <= 9'b11000111;
				8'b1001111: c <= 9'b10010;
				8'b1100101: c <= 9'b110111000;
				8'b1111110: c <= 9'b111101100;
				8'b1111100: c <= 9'b110111100;
				8'b1010110: c <= 9'b101011010;
				8'b110010: c <= 9'b1111000;
				8'b1101101: c <= 9'b110000111;
				8'b100011: c <= 9'b10001000;
				8'b1110101: c <= 9'b101000111;
				8'b1111101: c <= 9'b11100110;
				8'b101001: c <= 9'b1000110;
				8'b1010010: c <= 9'b10001101;
				8'b1011000: c <= 9'b10101011;
				8'b101110: c <= 9'b11111;
				8'b1000001: c <= 9'b101110011;
				default: c <= 9'b0;
			endcase
			9'b101111100 : case(di)
				8'b1000011: c <= 9'b11110010;
				8'b101000: c <= 9'b1100100;
				8'b111010: c <= 9'b10011011;
				8'b110110: c <= 9'b10001100;
				8'b1100100: c <= 9'b10000001;
				8'b1000000: c <= 9'b110101101;
				8'b1110110: c <= 9'b101011101;
				8'b100101: c <= 9'b101100110;
				8'b101111: c <= 9'b1111110;
				8'b100110: c <= 9'b111100100;
				8'b1100011: c <= 9'b110110110;
				8'b1001000: c <= 9'b10001010;
				8'b111000: c <= 9'b1111101;
				8'b110001: c <= 9'b1001011;
				8'b1010111: c <= 9'b100011111;
				8'b1001110: c <= 9'b1101010;
				8'b1101010: c <= 9'b11010100;
				8'b1001001: c <= 9'b1101;
				8'b1100000: c <= 9'b110010110;
				8'b110111: c <= 9'b111011111;
				8'b1011101: c <= 9'b10001011;
				8'b1011011: c <= 9'b10100011;
				8'b111001: c <= 9'b100101110;
				8'b1001010: c <= 9'b101010110;
				8'b110011: c <= 9'b10011010;
				8'b1101100: c <= 9'b101010100;
				8'b1110111: c <= 9'b10010011;
				8'b101011: c <= 9'b10010110;
				8'b1101011: c <= 9'b100100001;
				8'b111100: c <= 9'b1101010;
				8'b1000111: c <= 9'b10001010;
				8'b1011111: c <= 9'b101001;
				8'b1110100: c <= 9'b1010001;
				8'b101101: c <= 9'b100101110;
				8'b1010011: c <= 9'b11001011;
				8'b1100001: c <= 9'b110000111;
				8'b110101: c <= 9'b10111010;
				8'b1000100: c <= 9'b110010110;
				8'b1010001: c <= 9'b11011101;
				8'b1010100: c <= 9'b110001000;
				8'b1100110: c <= 9'b110100101;
				8'b101010: c <= 9'b10101010;
				8'b1011110: c <= 9'b11111110;
				8'b1100111: c <= 9'b10010110;
				8'b1011010: c <= 9'b100010000;
				8'b1000010: c <= 9'b110110;
				8'b111101: c <= 9'b11010111;
				8'b110000: c <= 9'b110110001;
				8'b111110: c <= 9'b1010001;
				8'b1100010: c <= 9'b111001111;
				8'b1110000: c <= 9'b1011011;
				8'b1101001: c <= 9'b11011110;
				8'b1110011: c <= 9'b10011000;
				8'b1001100: c <= 9'b11000011;
				8'b100001: c <= 9'b1110;
				8'b1000110: c <= 9'b10010100;
				8'b1110010: c <= 9'b111100000;
				8'b1010000: c <= 9'b100010010;
				8'b1111010: c <= 9'b101100010;
				8'b1010101: c <= 9'b100101100;
				8'b111011: c <= 9'b110110000;
				8'b1001101: c <= 9'b110111;
				8'b111111: c <= 9'b101000011;
				8'b1101110: c <= 9'b11110111;
				8'b1111011: c <= 9'b10111111;
				8'b1001011: c <= 9'b100010;
				8'b1101111: c <= 9'b110110;
				8'b1101000: c <= 9'b10100100;
				8'b101100: c <= 9'b111111000;
				8'b100100: c <= 9'b101101111;
				8'b1111000: c <= 9'b101111111;
				8'b1000101: c <= 9'b1101110;
				8'b1011001: c <= 9'b110011110;
				8'b110100: c <= 9'b111111000;
				8'b1111001: c <= 9'b11000011;
				8'b1110001: c <= 9'b1001101;
				8'b1001111: c <= 9'b11000010;
				8'b1100101: c <= 9'b10010;
				8'b1111110: c <= 9'b1100011;
				8'b1111100: c <= 9'b10010100;
				8'b1010110: c <= 9'b110100100;
				8'b110010: c <= 9'b111011110;
				8'b1101101: c <= 9'b100111111;
				8'b100011: c <= 9'b1000010;
				8'b1110101: c <= 9'b11110100;
				8'b1111101: c <= 9'b100110100;
				8'b101001: c <= 9'b111110101;
				8'b1010010: c <= 9'b100101;
				8'b1011000: c <= 9'b110100000;
				8'b101110: c <= 9'b111000000;
				8'b1000001: c <= 9'b11110000;
				default: c <= 9'b0;
			endcase
			9'b110110001 : case(di)
				8'b1000011: c <= 9'b100100;
				8'b101000: c <= 9'b110110011;
				8'b111010: c <= 9'b101001100;
				8'b110110: c <= 9'b101001000;
				8'b1100100: c <= 9'b11100111;
				8'b1000000: c <= 9'b101011;
				8'b1110110: c <= 9'b11110100;
				8'b100101: c <= 9'b11100111;
				8'b101111: c <= 9'b11010010;
				8'b100110: c <= 9'b110000001;
				8'b1100011: c <= 9'b111111110;
				8'b1001000: c <= 9'b100101011;
				8'b111000: c <= 9'b100110011;
				8'b110001: c <= 9'b10100101;
				8'b1010111: c <= 9'b110001110;
				8'b1001110: c <= 9'b100001011;
				8'b1101010: c <= 9'b110011001;
				8'b1001001: c <= 9'b110000011;
				8'b1100000: c <= 9'b111110101;
				8'b110111: c <= 9'b1110011;
				8'b1011101: c <= 9'b111000100;
				8'b1011011: c <= 9'b101111111;
				8'b111001: c <= 9'b110100110;
				8'b1001010: c <= 9'b11110110;
				8'b110011: c <= 9'b10110110;
				8'b1101100: c <= 9'b110110111;
				8'b1110111: c <= 9'b11101111;
				8'b101011: c <= 9'b100100000;
				8'b1101011: c <= 9'b10010101;
				8'b111100: c <= 9'b11100;
				8'b1000111: c <= 9'b100001100;
				8'b1011111: c <= 9'b101100011;
				8'b1110100: c <= 9'b100100001;
				8'b101101: c <= 9'b1010010;
				8'b1010011: c <= 9'b110111;
				8'b1100001: c <= 9'b10000010;
				8'b110101: c <= 9'b10101010;
				8'b1000100: c <= 9'b11011100;
				8'b1010001: c <= 9'b110000010;
				8'b1010100: c <= 9'b110100010;
				8'b1100110: c <= 9'b10100110;
				8'b101010: c <= 9'b100100011;
				8'b1011110: c <= 9'b111111101;
				8'b1100111: c <= 9'b111000101;
				8'b1011010: c <= 9'b110011100;
				8'b1000010: c <= 9'b110000111;
				8'b111101: c <= 9'b111011010;
				8'b110000: c <= 9'b11100;
				8'b111110: c <= 9'b1100010;
				8'b1100010: c <= 9'b1101000;
				8'b1110000: c <= 9'b10000;
				8'b1101001: c <= 9'b10100100;
				8'b1110011: c <= 9'b111111110;
				8'b1001100: c <= 9'b1101000;
				8'b100001: c <= 9'b1100001;
				8'b1000110: c <= 9'b101;
				8'b1110010: c <= 9'b1000000;
				8'b1010000: c <= 9'b1001011;
				8'b1111010: c <= 9'b110110000;
				8'b1010101: c <= 9'b111100111;
				8'b111011: c <= 9'b10010100;
				8'b1001101: c <= 9'b110110100;
				8'b111111: c <= 9'b101101011;
				8'b1101110: c <= 9'b111010100;
				8'b1111011: c <= 9'b100000101;
				8'b1001011: c <= 9'b100010010;
				8'b1101111: c <= 9'b10100000;
				8'b1101000: c <= 9'b111110110;
				8'b101100: c <= 9'b100111101;
				8'b100100: c <= 9'b111110000;
				8'b1111000: c <= 9'b111000101;
				8'b1000101: c <= 9'b100111010;
				8'b1011001: c <= 9'b110110011;
				8'b110100: c <= 9'b1000001;
				8'b1111001: c <= 9'b1101101;
				8'b1110001: c <= 9'b1110010;
				8'b1001111: c <= 9'b1011000;
				8'b1100101: c <= 9'b100010110;
				8'b1111110: c <= 9'b10100110;
				8'b1111100: c <= 9'b110010;
				8'b1010110: c <= 9'b110100100;
				8'b110010: c <= 9'b1000000;
				8'b1101101: c <= 9'b10101010;
				8'b100011: c <= 9'b1110111;
				8'b1110101: c <= 9'b11101010;
				8'b1111101: c <= 9'b11011010;
				8'b101001: c <= 9'b11110011;
				8'b1010010: c <= 9'b100110101;
				8'b1011000: c <= 9'b111011;
				8'b101110: c <= 9'b10110010;
				8'b1000001: c <= 9'b1111101;
				default: c <= 9'b0;
			endcase
			9'b11101010 : case(di)
				8'b1000011: c <= 9'b101001011;
				8'b101000: c <= 9'b10001101;
				8'b111010: c <= 9'b111001100;
				8'b110110: c <= 9'b110111011;
				8'b1100100: c <= 9'b11000001;
				8'b1000000: c <= 9'b111010111;
				8'b1110110: c <= 9'b111011111;
				8'b100101: c <= 9'b11110000;
				8'b101111: c <= 9'b10100101;
				8'b100110: c <= 9'b110011101;
				8'b1100011: c <= 9'b1101111;
				8'b1001000: c <= 9'b1010101;
				8'b111000: c <= 9'b101100011;
				8'b110001: c <= 9'b11100010;
				8'b1010111: c <= 9'b11100110;
				8'b1001110: c <= 9'b110100111;
				8'b1101010: c <= 9'b1100011;
				8'b1001001: c <= 9'b100101;
				8'b1100000: c <= 9'b10000001;
				8'b110111: c <= 9'b110010011;
				8'b1011101: c <= 9'b100;
				8'b1011011: c <= 9'b11001100;
				8'b111001: c <= 9'b100101100;
				8'b1001010: c <= 9'b101101011;
				8'b110011: c <= 9'b11111011;
				8'b1101100: c <= 9'b111100100;
				8'b1110111: c <= 9'b111000000;
				8'b101011: c <= 9'b1010000;
				8'b1101011: c <= 9'b1101010;
				8'b111100: c <= 9'b101001100;
				8'b1000111: c <= 9'b11;
				8'b1011111: c <= 9'b1010100;
				8'b1110100: c <= 9'b10011111;
				8'b101101: c <= 9'b1100111;
				8'b1010011: c <= 9'b111110011;
				8'b1100001: c <= 9'b100000101;
				8'b110101: c <= 9'b100101100;
				8'b1000100: c <= 9'b110011;
				8'b1010001: c <= 9'b111101100;
				8'b1010100: c <= 9'b111100101;
				8'b1100110: c <= 9'b11010001;
				8'b101010: c <= 9'b11101011;
				8'b1011110: c <= 9'b111001010;
				8'b1100111: c <= 9'b1001000;
				8'b1011010: c <= 9'b100000111;
				8'b1000010: c <= 9'b1000010;
				8'b111101: c <= 9'b111000010;
				8'b110000: c <= 9'b11100010;
				8'b111110: c <= 9'b11001101;
				8'b1100010: c <= 9'b100100111;
				8'b1110000: c <= 9'b110110000;
				8'b1101001: c <= 9'b111101101;
				8'b1110011: c <= 9'b101110010;
				8'b1001100: c <= 9'b110011110;
				8'b100001: c <= 9'b110010111;
				8'b1000110: c <= 9'b100001001;
				8'b1110010: c <= 9'b1000110;
				8'b1010000: c <= 9'b110111010;
				8'b1111010: c <= 9'b1001111;
				8'b1010101: c <= 9'b101010110;
				8'b111011: c <= 9'b1011010;
				8'b1001101: c <= 9'b100101010;
				8'b111111: c <= 9'b101111000;
				8'b1101110: c <= 9'b111001100;
				8'b1111011: c <= 9'b101100110;
				8'b1001011: c <= 9'b1111100;
				8'b1101111: c <= 9'b111101101;
				8'b1101000: c <= 9'b101110110;
				8'b101100: c <= 9'b100011000;
				8'b100100: c <= 9'b101000001;
				8'b1111000: c <= 9'b100001100;
				8'b1000101: c <= 9'b101000100;
				8'b1011001: c <= 9'b100001010;
				8'b110100: c <= 9'b1000010;
				8'b1111001: c <= 9'b10001011;
				8'b1110001: c <= 9'b111100101;
				8'b1001111: c <= 9'b100001;
				8'b1100101: c <= 9'b1011110;
				8'b1111110: c <= 9'b100101010;
				8'b1111100: c <= 9'b100100000;
				8'b1010110: c <= 9'b100000001;
				8'b110010: c <= 9'b1101100;
				8'b1101101: c <= 9'b1101001;
				8'b100011: c <= 9'b11010100;
				8'b1110101: c <= 9'b101101011;
				8'b1111101: c <= 9'b110000000;
				8'b101001: c <= 9'b11001001;
				8'b1010010: c <= 9'b1011100;
				8'b1011000: c <= 9'b1111101;
				8'b101110: c <= 9'b110111001;
				8'b1000001: c <= 9'b110110010;
				default: c <= 9'b0;
			endcase
			9'b1010100 : case(di)
				8'b1000011: c <= 9'b110100;
				8'b101000: c <= 9'b101100111;
				8'b111010: c <= 9'b11000110;
				8'b110110: c <= 9'b110100111;
				8'b1100100: c <= 9'b1001110;
				8'b1000000: c <= 9'b10001101;
				8'b1110110: c <= 9'b11010000;
				8'b100101: c <= 9'b111100010;
				8'b101111: c <= 9'b110111100;
				8'b100110: c <= 9'b110111110;
				8'b1100011: c <= 9'b110010;
				8'b1001000: c <= 9'b101000110;
				8'b111000: c <= 9'b10111111;
				8'b110001: c <= 9'b10010011;
				8'b1010111: c <= 9'b11001011;
				8'b1001110: c <= 9'b100011010;
				8'b1101010: c <= 9'b110001110;
				8'b1001001: c <= 9'b100011000;
				8'b1100000: c <= 9'b11010;
				8'b110111: c <= 9'b110110100;
				8'b1011101: c <= 9'b101010111;
				8'b1011011: c <= 9'b10111111;
				8'b111001: c <= 9'b100110000;
				8'b1001010: c <= 9'b1101000;
				8'b110011: c <= 9'b1010110;
				8'b1101100: c <= 9'b101000;
				8'b1110111: c <= 9'b1010111;
				8'b101011: c <= 9'b100000000;
				8'b1101011: c <= 9'b1000110;
				8'b111100: c <= 9'b101110010;
				8'b1000111: c <= 9'b110000001;
				8'b1011111: c <= 9'b100111101;
				8'b1110100: c <= 9'b100011;
				8'b101101: c <= 9'b100001;
				8'b1010011: c <= 9'b1110100;
				8'b1100001: c <= 9'b100000110;
				8'b110101: c <= 9'b11010011;
				8'b1000100: c <= 9'b100010100;
				8'b1010001: c <= 9'b101111110;
				8'b1010100: c <= 9'b100011010;
				8'b1100110: c <= 9'b111011011;
				8'b101010: c <= 9'b111101111;
				8'b1011110: c <= 9'b1011011;
				8'b1100111: c <= 9'b11000;
				8'b1011010: c <= 9'b10100010;
				8'b1000010: c <= 9'b11101111;
				8'b111101: c <= 9'b100011100;
				8'b110000: c <= 9'b100001010;
				8'b111110: c <= 9'b111011001;
				8'b1100010: c <= 9'b1011000;
				8'b1110000: c <= 9'b1011;
				8'b1101001: c <= 9'b100010100;
				8'b1110011: c <= 9'b110001010;
				8'b1001100: c <= 9'b1001000;
				8'b100001: c <= 9'b110100010;
				8'b1000110: c <= 9'b111111001;
				8'b1110010: c <= 9'b11;
				8'b1010000: c <= 9'b101111000;
				8'b1111010: c <= 9'b111101001;
				8'b1010101: c <= 9'b11100001;
				8'b111011: c <= 9'b100111;
				8'b1001101: c <= 9'b101011010;
				8'b111111: c <= 9'b111111010;
				8'b1101110: c <= 9'b1101101;
				8'b1111011: c <= 9'b101101011;
				8'b1001011: c <= 9'b100111110;
				8'b1101111: c <= 9'b1100000;
				8'b1101000: c <= 9'b100011000;
				8'b101100: c <= 9'b10100000;
				8'b100100: c <= 9'b11000011;
				8'b1111000: c <= 9'b10110;
				8'b1000101: c <= 9'b11000;
				8'b1011001: c <= 9'b1100101;
				8'b110100: c <= 9'b11001;
				8'b1111001: c <= 9'b110101;
				8'b1110001: c <= 9'b1001011;
				8'b1001111: c <= 9'b110111011;
				8'b1100101: c <= 9'b1100101;
				8'b1111110: c <= 9'b1100011;
				8'b1111100: c <= 9'b10101011;
				8'b1010110: c <= 9'b10111111;
				8'b110010: c <= 9'b100100011;
				8'b1101101: c <= 9'b10001010;
				8'b100011: c <= 9'b110110011;
				8'b1110101: c <= 9'b110111101;
				8'b1111101: c <= 9'b101100101;
				8'b101001: c <= 9'b1000;
				8'b1010010: c <= 9'b110100010;
				8'b1011000: c <= 9'b101001100;
				8'b101110: c <= 9'b10100010;
				8'b1000001: c <= 9'b111100010;
				default: c <= 9'b0;
			endcase
			9'b110111101 : case(di)
				8'b1000011: c <= 9'b110010;
				8'b101000: c <= 9'b110011110;
				8'b111010: c <= 9'b110110011;
				8'b110110: c <= 9'b1110100;
				8'b1100100: c <= 9'b110000011;
				8'b1000000: c <= 9'b11101111;
				8'b1110110: c <= 9'b1001110;
				8'b100101: c <= 9'b111100;
				8'b101111: c <= 9'b11011101;
				8'b100110: c <= 9'b111000111;
				8'b1100011: c <= 9'b1101001;
				8'b1001000: c <= 9'b100000001;
				8'b111000: c <= 9'b111010;
				8'b110001: c <= 9'b10010101;
				8'b1010111: c <= 9'b10011010;
				8'b1001110: c <= 9'b111101111;
				8'b1101010: c <= 9'b10011001;
				8'b1001001: c <= 9'b111011110;
				8'b1100000: c <= 9'b101100111;
				8'b110111: c <= 9'b100111101;
				8'b1011101: c <= 9'b101111001;
				8'b1011011: c <= 9'b1001011;
				8'b111001: c <= 9'b100011111;
				8'b1001010: c <= 9'b10000;
				8'b110011: c <= 9'b101110110;
				8'b1101100: c <= 9'b1001001;
				8'b1110111: c <= 9'b100000101;
				8'b101011: c <= 9'b100000111;
				8'b1101011: c <= 9'b10000001;
				8'b111100: c <= 9'b11011010;
				8'b1000111: c <= 9'b101011101;
				8'b1011111: c <= 9'b1011;
				8'b1110100: c <= 9'b10000001;
				8'b101101: c <= 9'b11100000;
				8'b1010011: c <= 9'b110010;
				8'b1100001: c <= 9'b101001000;
				8'b110101: c <= 9'b100010101;
				8'b1000100: c <= 9'b101010100;
				8'b1010001: c <= 9'b111111011;
				8'b1010100: c <= 9'b110110000;
				8'b1100110: c <= 9'b110010011;
				8'b101010: c <= 9'b11001111;
				8'b1011110: c <= 9'b10001001;
				8'b1100111: c <= 9'b101100100;
				8'b1011010: c <= 9'b10101011;
				8'b1000010: c <= 9'b11011000;
				8'b111101: c <= 9'b110000001;
				8'b110000: c <= 9'b1110001;
				8'b111110: c <= 9'b101010;
				8'b1100010: c <= 9'b11101001;
				8'b1110000: c <= 9'b111000000;
				8'b1101001: c <= 9'b101001001;
				8'b1110011: c <= 9'b1010;
				8'b1001100: c <= 9'b101000001;
				8'b100001: c <= 9'b101011110;
				8'b1000110: c <= 9'b100000111;
				8'b1110010: c <= 9'b100001101;
				8'b1010000: c <= 9'b101110110;
				8'b1111010: c <= 9'b11110101;
				8'b1010101: c <= 9'b1101101;
				8'b111011: c <= 9'b111011011;
				8'b1001101: c <= 9'b11000111;
				8'b111111: c <= 9'b1111001;
				8'b1101110: c <= 9'b11111000;
				8'b1111011: c <= 9'b10111001;
				8'b1001011: c <= 9'b111001000;
				8'b1101111: c <= 9'b11111;
				8'b1101000: c <= 9'b101010000;
				8'b101100: c <= 9'b10011;
				8'b100100: c <= 9'b110011100;
				8'b1111000: c <= 9'b111000000;
				8'b1000101: c <= 9'b111011100;
				8'b1011001: c <= 9'b10010110;
				8'b110100: c <= 9'b10011001;
				8'b1111001: c <= 9'b11001111;
				8'b1110001: c <= 9'b110000111;
				8'b1001111: c <= 9'b1011010;
				8'b1100101: c <= 9'b100010111;
				8'b1111110: c <= 9'b1011111;
				8'b1111100: c <= 9'b1001111;
				8'b1010110: c <= 9'b111110101;
				8'b110010: c <= 9'b100111001;
				8'b1101101: c <= 9'b11001111;
				8'b100011: c <= 9'b100010001;
				8'b1110101: c <= 9'b10100100;
				8'b1111101: c <= 9'b110111011;
				8'b101001: c <= 9'b101011;
				8'b1010010: c <= 9'b100100011;
				8'b1011000: c <= 9'b100010011;
				8'b101110: c <= 9'b1100010;
				8'b1000001: c <= 9'b101101111;
				default: c <= 9'b0;
			endcase
			9'b1010 : case(di)
				8'b1000011: c <= 9'b1000100;
				8'b101000: c <= 9'b110001010;
				8'b111010: c <= 9'b11010100;
				8'b110110: c <= 9'b110011111;
				8'b1100100: c <= 9'b110000010;
				8'b1000000: c <= 9'b100;
				8'b1110110: c <= 9'b101111010;
				8'b100101: c <= 9'b11000000;
				8'b101111: c <= 9'b100110000;
				8'b100110: c <= 9'b1010111;
				8'b1100011: c <= 9'b110000011;
				8'b1001000: c <= 9'b111001110;
				8'b111000: c <= 9'b110011100;
				8'b110001: c <= 9'b101111111;
				8'b1010111: c <= 9'b110011110;
				8'b1001110: c <= 9'b101001011;
				8'b1101010: c <= 9'b11000;
				8'b1001001: c <= 9'b110010110;
				8'b1100000: c <= 9'b11110011;
				8'b110111: c <= 9'b11101001;
				8'b1011101: c <= 9'b110100100;
				8'b1011011: c <= 9'b101100101;
				8'b111001: c <= 9'b110011001;
				8'b1001010: c <= 9'b11110100;
				8'b110011: c <= 9'b10110000;
				8'b1101100: c <= 9'b110101110;
				8'b1110111: c <= 9'b1011001;
				8'b101011: c <= 9'b111000110;
				8'b1101011: c <= 9'b100011001;
				8'b111100: c <= 9'b1000011;
				8'b1000111: c <= 9'b10010101;
				8'b1011111: c <= 9'b110110100;
				8'b1110100: c <= 9'b110010011;
				8'b101101: c <= 9'b11100100;
				8'b1010011: c <= 9'b1010011;
				8'b1100001: c <= 9'b110011010;
				8'b110101: c <= 9'b1010001;
				8'b1000100: c <= 9'b100101100;
				8'b1010001: c <= 9'b111111010;
				8'b1010100: c <= 9'b11110010;
				8'b1100110: c <= 9'b10100;
				8'b101010: c <= 9'b10100;
				8'b1011110: c <= 9'b1001110;
				8'b1100111: c <= 9'b110010011;
				8'b1011010: c <= 9'b10110110;
				8'b1000010: c <= 9'b1000000;
				8'b111101: c <= 9'b100010011;
				8'b110000: c <= 9'b111000110;
				8'b111110: c <= 9'b101110010;
				8'b1100010: c <= 9'b111111111;
				8'b1110000: c <= 9'b1000100;
				8'b1101001: c <= 9'b101101000;
				8'b1110011: c <= 9'b101100100;
				8'b1001100: c <= 9'b100110000;
				8'b100001: c <= 9'b100001011;
				8'b1000110: c <= 9'b100000101;
				8'b1110010: c <= 9'b1100101;
				8'b1010000: c <= 9'b11111000;
				8'b1111010: c <= 9'b110010110;
				8'b1010101: c <= 9'b110111;
				8'b111011: c <= 9'b11110110;
				8'b1001101: c <= 9'b100111010;
				8'b111111: c <= 9'b111111101;
				8'b1101110: c <= 9'b11110;
				8'b1111011: c <= 9'b100110010;
				8'b1001011: c <= 9'b1101110;
				8'b1101111: c <= 9'b110101;
				8'b1101000: c <= 9'b100011111;
				8'b101100: c <= 9'b10001011;
				8'b100100: c <= 9'b11101100;
				8'b1111000: c <= 9'b110111111;
				8'b1000101: c <= 9'b1111100;
				8'b1011001: c <= 9'b11111100;
				8'b110100: c <= 9'b11001110;
				8'b1111001: c <= 9'b101101;
				8'b1110001: c <= 9'b101010000;
				8'b1001111: c <= 9'b101100011;
				8'b1100101: c <= 9'b1110011;
				8'b1111110: c <= 9'b111101000;
				8'b1111100: c <= 9'b11000001;
				8'b1010110: c <= 9'b110001000;
				8'b110010: c <= 9'b111011100;
				8'b1101101: c <= 9'b111001001;
				8'b100011: c <= 9'b10000110;
				8'b1110101: c <= 9'b1001011;
				8'b1111101: c <= 9'b100101010;
				8'b101001: c <= 9'b110100001;
				8'b1010010: c <= 9'b100000100;
				8'b1011000: c <= 9'b111110001;
				8'b101110: c <= 9'b1000;
				8'b1000001: c <= 9'b111111110;
				default: c <= 9'b0;
			endcase
			9'b10110000 : case(di)
				8'b1000011: c <= 9'b11111;
				8'b101000: c <= 9'b11101101;
				8'b111010: c <= 9'b100010101;
				8'b110110: c <= 9'b110001101;
				8'b1100100: c <= 9'b101000000;
				8'b1000000: c <= 9'b101111000;
				8'b1110110: c <= 9'b10101000;
				8'b100101: c <= 9'b111010100;
				8'b101111: c <= 9'b11100000;
				8'b100110: c <= 9'b10010111;
				8'b1100011: c <= 9'b100111000;
				8'b1001000: c <= 9'b100001011;
				8'b111000: c <= 9'b100110110;
				8'b110001: c <= 9'b10011111;
				8'b1010111: c <= 9'b11111010;
				8'b1001110: c <= 9'b101110001;
				8'b1101010: c <= 9'b1000011;
				8'b1001001: c <= 9'b100010010;
				8'b1100000: c <= 9'b11010100;
				8'b110111: c <= 9'b101011111;
				8'b1011101: c <= 9'b1110111;
				8'b1011011: c <= 9'b101100;
				8'b111001: c <= 9'b101100101;
				8'b1001010: c <= 9'b100001001;
				8'b110011: c <= 9'b101101110;
				8'b1101100: c <= 9'b100100000;
				8'b1110111: c <= 9'b1000110;
				8'b101011: c <= 9'b11101100;
				8'b1101011: c <= 9'b100001111;
				8'b111100: c <= 9'b110101101;
				8'b1000111: c <= 9'b110110010;
				8'b1011111: c <= 9'b11001011;
				8'b1110100: c <= 9'b101101010;
				8'b101101: c <= 9'b1011011;
				8'b1010011: c <= 9'b100000111;
				8'b1100001: c <= 9'b110111000;
				8'b110101: c <= 9'b101111000;
				8'b1000100: c <= 9'b110101101;
				8'b1010001: c <= 9'b110110011;
				8'b1010100: c <= 9'b110111010;
				8'b1100110: c <= 9'b110011010;
				8'b101010: c <= 9'b1010110;
				8'b1011110: c <= 9'b111001100;
				8'b1100111: c <= 9'b10101111;
				8'b1011010: c <= 9'b111111010;
				8'b1000010: c <= 9'b101000;
				8'b111101: c <= 9'b10010101;
				8'b110000: c <= 9'b10001110;
				8'b111110: c <= 9'b100001010;
				8'b1100010: c <= 9'b100111;
				8'b1110000: c <= 9'b11110011;
				8'b1101001: c <= 9'b111001001;
				8'b1110011: c <= 9'b1101100;
				8'b1001100: c <= 9'b110011011;
				8'b100001: c <= 9'b101110111;
				8'b1000110: c <= 9'b11110101;
				8'b1110010: c <= 9'b100111000;
				8'b1010000: c <= 9'b111010100;
				8'b1111010: c <= 9'b1110011;
				8'b1010101: c <= 9'b110100000;
				8'b111011: c <= 9'b11111010;
				8'b1001101: c <= 9'b11100011;
				8'b111111: c <= 9'b110100011;
				8'b1101110: c <= 9'b11111000;
				8'b1111011: c <= 9'b110110110;
				8'b1001011: c <= 9'b111001010;
				8'b1101111: c <= 9'b100101111;
				8'b1101000: c <= 9'b110101111;
				8'b101100: c <= 9'b111110110;
				8'b100100: c <= 9'b1000001;
				8'b1111000: c <= 9'b110011011;
				8'b1000101: c <= 9'b111001001;
				8'b1011001: c <= 9'b101110110;
				8'b110100: c <= 9'b110111;
				8'b1111001: c <= 9'b1010111;
				8'b1110001: c <= 9'b101000111;
				8'b1001111: c <= 9'b10100101;
				8'b1100101: c <= 9'b110010;
				8'b1111110: c <= 9'b111101101;
				8'b1111100: c <= 9'b110110110;
				8'b1010110: c <= 9'b100100000;
				8'b110010: c <= 9'b101010100;
				8'b1101101: c <= 9'b10100101;
				8'b100011: c <= 9'b110010001;
				8'b1110101: c <= 9'b11110011;
				8'b1111101: c <= 9'b1000111;
				8'b101001: c <= 9'b1100;
				8'b1010010: c <= 9'b10100;
				8'b1011000: c <= 9'b110010011;
				8'b101110: c <= 9'b1101001;
				8'b1000001: c <= 9'b1111011;
				default: c <= 9'b0;
			endcase
			9'b101000000 : case(di)
				8'b1000011: c <= 9'b110100;
				8'b101000: c <= 9'b100111;
				8'b111010: c <= 9'b100100111;
				8'b110110: c <= 9'b101110;
				8'b1100100: c <= 9'b11000010;
				8'b1000000: c <= 9'b101001000;
				8'b1110110: c <= 9'b111011100;
				8'b100101: c <= 9'b11101111;
				8'b101111: c <= 9'b101100111;
				8'b100110: c <= 9'b101110010;
				8'b1100011: c <= 9'b101001010;
				8'b1001000: c <= 9'b1000111;
				8'b111000: c <= 9'b11010011;
				8'b110001: c <= 9'b11101011;
				8'b1010111: c <= 9'b1001001;
				8'b1001110: c <= 9'b10010;
				8'b1101010: c <= 9'b1010111;
				8'b1001001: c <= 9'b10001101;
				8'b1100000: c <= 9'b100000011;
				8'b110111: c <= 9'b11001111;
				8'b1011101: c <= 9'b10111100;
				8'b1011011: c <= 9'b10111110;
				8'b111001: c <= 9'b101110111;
				8'b1001010: c <= 9'b1011001;
				8'b110011: c <= 9'b101010111;
				8'b1101100: c <= 9'b1111010;
				8'b1110111: c <= 9'b1011010;
				8'b101011: c <= 9'b101101011;
				8'b1101011: c <= 9'b110001000;
				8'b111100: c <= 9'b110011011;
				8'b1000111: c <= 9'b101010011;
				8'b1011111: c <= 9'b111110111;
				8'b1110100: c <= 9'b110010010;
				8'b101101: c <= 9'b110010011;
				8'b1010011: c <= 9'b110110110;
				8'b1100001: c <= 9'b111100;
				8'b110101: c <= 9'b100001011;
				8'b1000100: c <= 9'b100010;
				8'b1010001: c <= 9'b1101110;
				8'b1010100: c <= 9'b1100;
				8'b1100110: c <= 9'b10011011;
				8'b101010: c <= 9'b111111110;
				8'b1011110: c <= 9'b1001011;
				8'b1100111: c <= 9'b11110;
				8'b1011010: c <= 9'b101101011;
				8'b1000010: c <= 9'b100111010;
				8'b111101: c <= 9'b10111011;
				8'b110000: c <= 9'b110101100;
				8'b111110: c <= 9'b11000110;
				8'b1100010: c <= 9'b11011;
				8'b1110000: c <= 9'b11011010;
				8'b1101001: c <= 9'b101101;
				8'b1110011: c <= 9'b110000001;
				8'b1001100: c <= 9'b10100110;
				8'b100001: c <= 9'b10010011;
				8'b1000110: c <= 9'b11101011;
				8'b1110010: c <= 9'b110011110;
				8'b1010000: c <= 9'b100100000;
				8'b1111010: c <= 9'b101011110;
				8'b1010101: c <= 9'b110010001;
				8'b111011: c <= 9'b110101111;
				8'b1001101: c <= 9'b111001110;
				8'b111111: c <= 9'b111100110;
				8'b1101110: c <= 9'b10111010;
				8'b1111011: c <= 9'b1110100;
				8'b1001011: c <= 9'b1101;
				8'b1101111: c <= 9'b1000001;
				8'b1101000: c <= 9'b101100011;
				8'b101100: c <= 9'b1100111;
				8'b100100: c <= 9'b101110001;
				8'b1111000: c <= 9'b101111010;
				8'b1000101: c <= 9'b101111010;
				8'b1011001: c <= 9'b1001110;
				8'b110100: c <= 9'b11011001;
				8'b1111001: c <= 9'b101100001;
				8'b1110001: c <= 9'b10100;
				8'b1001111: c <= 9'b110000;
				8'b1100101: c <= 9'b10101011;
				8'b1111110: c <= 9'b1011010;
				8'b1111100: c <= 9'b111101010;
				8'b1010110: c <= 9'b1000100;
				8'b110010: c <= 9'b1100100;
				8'b1101101: c <= 9'b111100110;
				8'b100011: c <= 9'b100001011;
				8'b1110101: c <= 9'b111010000;
				8'b1111101: c <= 9'b101001111;
				8'b101001: c <= 9'b101110;
				8'b1010010: c <= 9'b10110010;
				8'b1011000: c <= 9'b100101001;
				8'b101110: c <= 9'b110111110;
				8'b1000001: c <= 9'b100011000;
				default: c <= 9'b0;
			endcase
			9'b111110111 : case(di)
				8'b1000011: c <= 9'b10100101;
				8'b101000: c <= 9'b111010110;
				8'b111010: c <= 9'b1100110;
				8'b110110: c <= 9'b111001001;
				8'b1100100: c <= 9'b11100101;
				8'b1000000: c <= 9'b11001;
				8'b1110110: c <= 9'b10010010;
				8'b100101: c <= 9'b11110001;
				8'b101111: c <= 9'b100100;
				8'b100110: c <= 9'b101011000;
				8'b1100011: c <= 9'b10110001;
				8'b1001000: c <= 9'b100001100;
				8'b111000: c <= 9'b1000;
				8'b110001: c <= 9'b11101011;
				8'b1010111: c <= 9'b111000000;
				8'b1001110: c <= 9'b111110110;
				8'b1101010: c <= 9'b100100010;
				8'b1001001: c <= 9'b1010000;
				8'b1100000: c <= 9'b101101110;
				8'b110111: c <= 9'b11011001;
				8'b1011101: c <= 9'b1001001;
				8'b1011011: c <= 9'b10011001;
				8'b111001: c <= 9'b111011010;
				8'b1001010: c <= 9'b1100;
				8'b110011: c <= 9'b10011001;
				8'b1101100: c <= 9'b110111000;
				8'b1110111: c <= 9'b11100100;
				8'b101011: c <= 9'b10011000;
				8'b1101011: c <= 9'b11110101;
				8'b111100: c <= 9'b110110010;
				8'b1000111: c <= 9'b11001000;
				8'b1011111: c <= 9'b100010010;
				8'b1110100: c <= 9'b1011000;
				8'b101101: c <= 9'b101010011;
				8'b1010011: c <= 9'b1011000;
				8'b1100001: c <= 9'b11010100;
				8'b110101: c <= 9'b11100010;
				8'b1000100: c <= 9'b1010001;
				8'b1010001: c <= 9'b10110;
				8'b1010100: c <= 9'b11001110;
				8'b1100110: c <= 9'b1101;
				8'b101010: c <= 9'b101001000;
				8'b1011110: c <= 9'b1010001;
				8'b1100111: c <= 9'b110010001;
				8'b1011010: c <= 9'b10111111;
				8'b1000010: c <= 9'b101010011;
				8'b111101: c <= 9'b111000000;
				8'b110000: c <= 9'b111100011;
				8'b111110: c <= 9'b100001001;
				8'b1100010: c <= 9'b100001010;
				8'b1110000: c <= 9'b11111011;
				8'b1101001: c <= 9'b101101010;
				8'b1110011: c <= 9'b101;
				8'b1001100: c <= 9'b111100110;
				8'b100001: c <= 9'b101101100;
				8'b1000110: c <= 9'b11000;
				8'b1110010: c <= 9'b10011010;
				8'b1010000: c <= 9'b10000;
				8'b1111010: c <= 9'b11110100;
				8'b1010101: c <= 9'b100101100;
				8'b111011: c <= 9'b100001001;
				8'b1001101: c <= 9'b11011001;
				8'b111111: c <= 9'b10100111;
				8'b1101110: c <= 9'b10101000;
				8'b1111011: c <= 9'b100111000;
				8'b1001011: c <= 9'b1101;
				8'b1101111: c <= 9'b111111;
				8'b1101000: c <= 9'b111111000;
				8'b101100: c <= 9'b11000110;
				8'b100100: c <= 9'b110000110;
				8'b1111000: c <= 9'b110001;
				8'b1000101: c <= 9'b100010101;
				8'b1011001: c <= 9'b11110101;
				8'b110100: c <= 9'b111100001;
				8'b1111001: c <= 9'b100010001;
				8'b1110001: c <= 9'b100001110;
				8'b1001111: c <= 9'b111000110;
				8'b1100101: c <= 9'b111010111;
				8'b1111110: c <= 9'b1001101;
				8'b1111100: c <= 9'b110000101;
				8'b1010110: c <= 9'b10110111;
				8'b110010: c <= 9'b100100010;
				8'b1101101: c <= 9'b101110110;
				8'b100011: c <= 9'b1111011;
				8'b1110101: c <= 9'b100101010;
				8'b1111101: c <= 9'b101100;
				8'b101001: c <= 9'b110011100;
				8'b1010010: c <= 9'b110010100;
				8'b1011000: c <= 9'b11000001;
				8'b101110: c <= 9'b101011000;
				8'b1000001: c <= 9'b10000011;
				default: c <= 9'b0;
			endcase
			9'b10010010 : case(di)
				8'b1000011: c <= 9'b101011111;
				8'b101000: c <= 9'b111100010;
				8'b111010: c <= 9'b111010;
				8'b110110: c <= 9'b1011001;
				8'b1100100: c <= 9'b1010011;
				8'b1000000: c <= 9'b1000111;
				8'b1110110: c <= 9'b110010011;
				8'b100101: c <= 9'b111111000;
				8'b101111: c <= 9'b10111111;
				8'b100110: c <= 9'b1010101;
				8'b1100011: c <= 9'b111101000;
				8'b1001000: c <= 9'b10110100;
				8'b111000: c <= 9'b110010011;
				8'b110001: c <= 9'b101010010;
				8'b1010111: c <= 9'b100101100;
				8'b1001110: c <= 9'b111001010;
				8'b1101010: c <= 9'b100100111;
				8'b1001001: c <= 9'b101010011;
				8'b1100000: c <= 9'b11001010;
				8'b110111: c <= 9'b1101001;
				8'b1011101: c <= 9'b110011011;
				8'b1011011: c <= 9'b11101100;
				8'b111001: c <= 9'b100110011;
				8'b1001010: c <= 9'b1000;
				8'b110011: c <= 9'b10001;
				8'b1101100: c <= 9'b10101101;
				8'b1110111: c <= 9'b11100111;
				8'b101011: c <= 9'b100001001;
				8'b1101011: c <= 9'b101100100;
				8'b111100: c <= 9'b11001001;
				8'b1000111: c <= 9'b101110001;
				8'b1011111: c <= 9'b101011010;
				8'b1110100: c <= 9'b101010111;
				8'b101101: c <= 9'b111001100;
				8'b1010011: c <= 9'b101100;
				8'b1100001: c <= 9'b101101110;
				8'b110101: c <= 9'b110011000;
				8'b1000100: c <= 9'b10100110;
				8'b1010001: c <= 9'b111101;
				8'b1010100: c <= 9'b111101111;
				8'b1100110: c <= 9'b1001101;
				8'b101010: c <= 9'b100001111;
				8'b1011110: c <= 9'b110110100;
				8'b1100111: c <= 9'b111000101;
				8'b1011010: c <= 9'b111010110;
				8'b1000010: c <= 9'b101100011;
				8'b111101: c <= 9'b1100;
				8'b110000: c <= 9'b11001110;
				8'b111110: c <= 9'b111001111;
				8'b1100010: c <= 9'b11100;
				8'b1110000: c <= 9'b10110;
				8'b1101001: c <= 9'b1111;
				8'b1110011: c <= 9'b10000101;
				8'b1001100: c <= 9'b11110001;
				8'b100001: c <= 9'b110011001;
				8'b1000110: c <= 9'b101010011;
				8'b1110010: c <= 9'b11111110;
				8'b1010000: c <= 9'b1101001;
				8'b1111010: c <= 9'b1001011;
				8'b1010101: c <= 9'b1111101;
				8'b111011: c <= 9'b110000001;
				8'b1001101: c <= 9'b111100101;
				8'b111111: c <= 9'b10111101;
				8'b1101110: c <= 9'b100111001;
				8'b1111011: c <= 9'b10001011;
				8'b1001011: c <= 9'b110111001;
				8'b1101111: c <= 9'b11110101;
				8'b1101000: c <= 9'b1101;
				8'b101100: c <= 9'b10110010;
				8'b100100: c <= 9'b11101011;
				8'b1111000: c <= 9'b101100;
				8'b1000101: c <= 9'b100010010;
				8'b1011001: c <= 9'b100011;
				8'b110100: c <= 9'b110100110;
				8'b1111001: c <= 9'b111001110;
				8'b1110001: c <= 9'b10001111;
				8'b1001111: c <= 9'b10000010;
				8'b1100101: c <= 9'b100100010;
				8'b1111110: c <= 9'b11001010;
				8'b1111100: c <= 9'b101110;
				8'b1010110: c <= 9'b101100101;
				8'b110010: c <= 9'b110100010;
				8'b1101101: c <= 9'b11100010;
				8'b100011: c <= 9'b101110101;
				8'b1110101: c <= 9'b111010010;
				8'b1111101: c <= 9'b110111000;
				8'b101001: c <= 9'b100101101;
				8'b1010010: c <= 9'b101100010;
				8'b1011000: c <= 9'b11111001;
				8'b101110: c <= 9'b100110000;
				8'b1000001: c <= 9'b11011;
				default: c <= 9'b0;
			endcase
			9'b10001 : case(di)
				8'b1000011: c <= 9'b1101;
				8'b101000: c <= 9'b101101;
				8'b111010: c <= 9'b110101101;
				8'b110110: c <= 9'b1000000;
				8'b1100100: c <= 9'b100010001;
				8'b1000000: c <= 9'b101110;
				8'b1110110: c <= 9'b1001110;
				8'b100101: c <= 9'b111110110;
				8'b101111: c <= 9'b10011010;
				8'b100110: c <= 9'b111000111;
				8'b1100011: c <= 9'b101001000;
				8'b1001000: c <= 9'b101;
				8'b111000: c <= 9'b1111001;
				8'b110001: c <= 9'b101011000;
				8'b1010111: c <= 9'b110011011;
				8'b1001110: c <= 9'b110011000;
				8'b1101010: c <= 9'b1010110;
				8'b1001001: c <= 9'b1001111;
				8'b1100000: c <= 9'b110000111;
				8'b110111: c <= 9'b100111011;
				8'b1011101: c <= 9'b100111110;
				8'b1011011: c <= 9'b100111011;
				8'b111001: c <= 9'b11110101;
				8'b1001010: c <= 9'b101100100;
				8'b110011: c <= 9'b101111111;
				8'b1101100: c <= 9'b11101;
				8'b1110111: c <= 9'b111001100;
				8'b101011: c <= 9'b111100000;
				8'b1101011: c <= 9'b100011;
				8'b111100: c <= 9'b111101000;
				8'b1000111: c <= 9'b11001;
				8'b1011111: c <= 9'b1001001;
				8'b1110100: c <= 9'b100011;
				8'b101101: c <= 9'b10101000;
				8'b1010011: c <= 9'b1100010;
				8'b1100001: c <= 9'b10100;
				8'b110101: c <= 9'b111011001;
				8'b1000100: c <= 9'b111111;
				8'b1010001: c <= 9'b111000;
				8'b1010100: c <= 9'b101011111;
				8'b1100110: c <= 9'b101100;
				8'b101010: c <= 9'b10011010;
				8'b1011110: c <= 9'b10101101;
				8'b1100111: c <= 9'b11011010;
				8'b1011010: c <= 9'b101010101;
				8'b1000010: c <= 9'b111010110;
				8'b111101: c <= 9'b10001001;
				8'b110000: c <= 9'b10100;
				8'b111110: c <= 9'b100000110;
				8'b1100010: c <= 9'b100111010;
				8'b1110000: c <= 9'b100110110;
				8'b1101001: c <= 9'b1111100;
				8'b1110011: c <= 9'b101101001;
				8'b1001100: c <= 9'b100011001;
				8'b100001: c <= 9'b10011001;
				8'b1000110: c <= 9'b1101;
				8'b1110010: c <= 9'b100000;
				8'b1010000: c <= 9'b11011110;
				8'b1111010: c <= 9'b111110110;
				8'b1010101: c <= 9'b1101010;
				8'b111011: c <= 9'b101001111;
				8'b1001101: c <= 9'b111000111;
				8'b111111: c <= 9'b11001110;
				8'b1101110: c <= 9'b101010110;
				8'b1111011: c <= 9'b1010001;
				8'b1001011: c <= 9'b101000110;
				8'b1101111: c <= 9'b111000000;
				8'b1101000: c <= 9'b10000101;
				8'b101100: c <= 9'b10110001;
				8'b100100: c <= 9'b1010111;
				8'b1111000: c <= 9'b111;
				8'b1000101: c <= 9'b101001011;
				8'b1011001: c <= 9'b10111010;
				8'b110100: c <= 9'b11000011;
				8'b1111001: c <= 9'b100101000;
				8'b1110001: c <= 9'b10010011;
				8'b1001111: c <= 9'b10111101;
				8'b1100101: c <= 9'b10000110;
				8'b1111110: c <= 9'b1100010;
				8'b1111100: c <= 9'b101100010;
				8'b1010110: c <= 9'b101101001;
				8'b110010: c <= 9'b10111000;
				8'b1101101: c <= 9'b100101;
				8'b100011: c <= 9'b1101110;
				8'b1110101: c <= 9'b101011;
				8'b1111101: c <= 9'b1010000;
				8'b101001: c <= 9'b110000000;
				8'b1010010: c <= 9'b1101;
				8'b1011000: c <= 9'b10111011;
				8'b101110: c <= 9'b1111;
				8'b1000001: c <= 9'b101000101;
				default: c <= 9'b0;
			endcase
			9'b100000 : case(di)
				8'b1000011: c <= 9'b1010001;
				8'b101000: c <= 9'b100000010;
				8'b111010: c <= 9'b100100110;
				8'b110110: c <= 9'b111010;
				8'b1100100: c <= 9'b110111011;
				8'b1000000: c <= 9'b10100100;
				8'b1110110: c <= 9'b110100100;
				8'b100101: c <= 9'b100110110;
				8'b101111: c <= 9'b101010011;
				8'b100110: c <= 9'b101100110;
				8'b1100011: c <= 9'b101010111;
				8'b1001000: c <= 9'b110001;
				8'b111000: c <= 9'b1110;
				8'b110001: c <= 9'b10100001;
				8'b1010111: c <= 9'b110101100;
				8'b1001110: c <= 9'b101110101;
				8'b1101010: c <= 9'b1110001;
				8'b1001001: c <= 9'b101101010;
				8'b1100000: c <= 9'b100010101;
				8'b110111: c <= 9'b101011;
				8'b1011101: c <= 9'b11000001;
				8'b1011011: c <= 9'b10001000;
				8'b111001: c <= 9'b111011001;
				8'b1001010: c <= 9'b100110010;
				8'b110011: c <= 9'b111100110;
				8'b1101100: c <= 9'b1000;
				8'b1110111: c <= 9'b1001010;
				8'b101011: c <= 9'b11101101;
				8'b1101011: c <= 9'b101100101;
				8'b111100: c <= 9'b100110110;
				8'b1000111: c <= 9'b101011110;
				8'b1011111: c <= 9'b110111111;
				8'b1110100: c <= 9'b100110000;
				8'b101101: c <= 9'b110001000;
				8'b1010011: c <= 9'b10010111;
				8'b1100001: c <= 9'b111001011;
				8'b110101: c <= 9'b10000101;
				8'b1000100: c <= 9'b110011011;
				8'b1010001: c <= 9'b110100010;
				8'b1010100: c <= 9'b11011;
				8'b1100110: c <= 9'b100001;
				8'b101010: c <= 9'b1011110;
				8'b1011110: c <= 9'b11111100;
				8'b1100111: c <= 9'b101011001;
				8'b1011010: c <= 9'b10111100;
				8'b1000010: c <= 9'b1011000;
				8'b111101: c <= 9'b100111001;
				8'b110000: c <= 9'b1100100;
				8'b111110: c <= 9'b1001011;
				8'b1100010: c <= 9'b10100000;
				8'b1110000: c <= 9'b111111110;
				8'b1101001: c <= 9'b111000101;
				8'b1110011: c <= 9'b11010100;
				8'b1001100: c <= 9'b1111110;
				8'b100001: c <= 9'b10011011;
				8'b1000110: c <= 9'b1111001;
				8'b1110010: c <= 9'b111100;
				8'b1010000: c <= 9'b101010100;
				8'b1111010: c <= 9'b10011001;
				8'b1010101: c <= 9'b101100000;
				8'b111011: c <= 9'b110110101;
				8'b1001101: c <= 9'b10001000;
				8'b111111: c <= 9'b1010110;
				8'b1101110: c <= 9'b100001;
				8'b1111011: c <= 9'b11011101;
				8'b1001011: c <= 9'b101011110;
				8'b1101111: c <= 9'b101101010;
				8'b1101000: c <= 9'b101100111;
				8'b101100: c <= 9'b1101000;
				8'b100100: c <= 9'b11010111;
				8'b1111000: c <= 9'b1011001;
				8'b1000101: c <= 9'b101010111;
				8'b1011001: c <= 9'b111111110;
				8'b110100: c <= 9'b1110000;
				8'b1111001: c <= 9'b11001101;
				8'b1110001: c <= 9'b10110110;
				8'b1001111: c <= 9'b11001110;
				8'b1100101: c <= 9'b100010100;
				8'b1111110: c <= 9'b111100100;
				8'b1111100: c <= 9'b100110;
				8'b1010110: c <= 9'b111101110;
				8'b110010: c <= 9'b110011011;
				8'b1101101: c <= 9'b1101101;
				8'b100011: c <= 9'b100000101;
				8'b1110101: c <= 9'b10010101;
				8'b1111101: c <= 9'b111001001;
				8'b101001: c <= 9'b110100011;
				8'b1010010: c <= 9'b100101010;
				8'b1011000: c <= 9'b1111101;
				8'b101110: c <= 9'b11000111;
				8'b1000001: c <= 9'b1101010;
				default: c <= 9'b0;
			endcase
			9'b10100001 : case(di)
				8'b1000011: c <= 9'b10000000;
				8'b101000: c <= 9'b1001000;
				8'b111010: c <= 9'b101111000;
				8'b110110: c <= 9'b10000;
				8'b1100100: c <= 9'b111011001;
				8'b1000000: c <= 9'b11001001;
				8'b1110110: c <= 9'b100100010;
				8'b100101: c <= 9'b11000001;
				8'b101111: c <= 9'b1010000;
				8'b100110: c <= 9'b100111001;
				8'b1100011: c <= 9'b1011010;
				8'b1001000: c <= 9'b111011110;
				8'b111000: c <= 9'b101100010;
				8'b110001: c <= 9'b101011101;
				8'b1010111: c <= 9'b111011010;
				8'b1001110: c <= 9'b10100110;
				8'b1101010: c <= 9'b1010110;
				8'b1001001: c <= 9'b10010101;
				8'b1100000: c <= 9'b1000011;
				8'b110111: c <= 9'b110010100;
				8'b1011101: c <= 9'b100100101;
				8'b1011011: c <= 9'b110111000;
				8'b111001: c <= 9'b10101110;
				8'b1001010: c <= 9'b100101000;
				8'b110011: c <= 9'b100001011;
				8'b1101100: c <= 9'b1111111;
				8'b1110111: c <= 9'b10111;
				8'b101011: c <= 9'b111111010;
				8'b1101011: c <= 9'b101011;
				8'b111100: c <= 9'b110101110;
				8'b1000111: c <= 9'b11010100;
				8'b1011111: c <= 9'b110111100;
				8'b1110100: c <= 9'b1000110;
				8'b101101: c <= 9'b1101110;
				8'b1010011: c <= 9'b110001000;
				8'b1100001: c <= 9'b100110011;
				8'b110101: c <= 9'b111001011;
				8'b1000100: c <= 9'b110011110;
				8'b1010001: c <= 9'b11100110;
				8'b1010100: c <= 9'b11110001;
				8'b1100110: c <= 9'b110110000;
				8'b101010: c <= 9'b100110000;
				8'b1011110: c <= 9'b110001110;
				8'b1100111: c <= 9'b1001100;
				8'b1011010: c <= 9'b100010101;
				8'b1000010: c <= 9'b101110111;
				8'b111101: c <= 9'b1011011;
				8'b110000: c <= 9'b100001111;
				8'b111110: c <= 9'b1111101;
				8'b1100010: c <= 9'b1101100;
				8'b1110000: c <= 9'b110101101;
				8'b1101001: c <= 9'b101010010;
				8'b1110011: c <= 9'b11110101;
				8'b1001100: c <= 9'b111011000;
				8'b100001: c <= 9'b1011111;
				8'b1000110: c <= 9'b10101000;
				8'b1110010: c <= 9'b10101001;
				8'b1010000: c <= 9'b111010010;
				8'b1111010: c <= 9'b100001001;
				8'b1010101: c <= 9'b101011110;
				8'b111011: c <= 9'b1101101;
				8'b1001101: c <= 9'b101101101;
				8'b111111: c <= 9'b11101;
				8'b1101110: c <= 9'b10101100;
				8'b1111011: c <= 9'b111101100;
				8'b1001011: c <= 9'b110110100;
				8'b1101111: c <= 9'b1010011;
				8'b1101000: c <= 9'b100011111;
				8'b101100: c <= 9'b100110101;
				8'b100100: c <= 9'b10101101;
				8'b1111000: c <= 9'b1010011;
				8'b1000101: c <= 9'b100010011;
				8'b1011001: c <= 9'b1000100;
				8'b110100: c <= 9'b1101110;
				8'b1111001: c <= 9'b101111001;
				8'b1110001: c <= 9'b111000000;
				8'b1001111: c <= 9'b11101100;
				8'b1100101: c <= 9'b100100110;
				8'b1111110: c <= 9'b101101100;
				8'b1111100: c <= 9'b111001110;
				8'b1010110: c <= 9'b111010;
				8'b110010: c <= 9'b1;
				8'b1101101: c <= 9'b111010000;
				8'b100011: c <= 9'b100001100;
				8'b1110101: c <= 9'b1000011;
				8'b1111101: c <= 9'b100010011;
				8'b101001: c <= 9'b100100001;
				8'b1010010: c <= 9'b11110011;
				8'b1011000: c <= 9'b10101010;
				8'b101110: c <= 9'b101101000;
				8'b1000001: c <= 9'b101010000;
				default: c <= 9'b0;
			endcase
			9'b111011000 : case(di)
				8'b1000011: c <= 9'b11001110;
				8'b101000: c <= 9'b11010100;
				8'b111010: c <= 9'b1011100;
				8'b110110: c <= 9'b11011100;
				8'b1100100: c <= 9'b1001001;
				8'b1000000: c <= 9'b110001110;
				8'b1110110: c <= 9'b100011101;
				8'b100101: c <= 9'b111001101;
				8'b101111: c <= 9'b100000011;
				8'b100110: c <= 9'b111100101;
				8'b1100011: c <= 9'b111000110;
				8'b1001000: c <= 9'b10111101;
				8'b111000: c <= 9'b10010101;
				8'b110001: c <= 9'b111000011;
				8'b1010111: c <= 9'b110100010;
				8'b1001110: c <= 9'b1;
				8'b1101010: c <= 9'b101011111;
				8'b1001001: c <= 9'b110010110;
				8'b1100000: c <= 9'b1110111;
				8'b110111: c <= 9'b1000000;
				8'b1011101: c <= 9'b111111;
				8'b1011011: c <= 9'b111111011;
				8'b111001: c <= 9'b111011;
				8'b1001010: c <= 9'b11000111;
				8'b110011: c <= 9'b101001000;
				8'b1101100: c <= 9'b11000;
				8'b1110111: c <= 9'b110100001;
				8'b101011: c <= 9'b10000111;
				8'b1101011: c <= 9'b111011100;
				8'b111100: c <= 9'b111100101;
				8'b1000111: c <= 9'b100100011;
				8'b1011111: c <= 9'b110101110;
				8'b1110100: c <= 9'b1000010;
				8'b101101: c <= 9'b1001101;
				8'b1010011: c <= 9'b110001000;
				8'b1100001: c <= 9'b110111001;
				8'b110101: c <= 9'b1001001;
				8'b1000100: c <= 9'b11011010;
				8'b1010001: c <= 9'b10100111;
				8'b1010100: c <= 9'b111000100;
				8'b1100110: c <= 9'b100001100;
				8'b101010: c <= 9'b111000101;
				8'b1011110: c <= 9'b110110100;
				8'b1100111: c <= 9'b101100110;
				8'b1011010: c <= 9'b110111;
				8'b1000010: c <= 9'b111001001;
				8'b111101: c <= 9'b111010001;
				8'b110000: c <= 9'b111111111;
				8'b111110: c <= 9'b11110001;
				8'b1100010: c <= 9'b100001111;
				8'b1110000: c <= 9'b11101000;
				8'b1101001: c <= 9'b110010011;
				8'b1110011: c <= 9'b11001011;
				8'b1001100: c <= 9'b1110111;
				8'b100001: c <= 9'b100100010;
				8'b1000110: c <= 9'b10010101;
				8'b1110010: c <= 9'b10010111;
				8'b1010000: c <= 9'b1011110;
				8'b1111010: c <= 9'b110110101;
				8'b1010101: c <= 9'b101110111;
				8'b111011: c <= 9'b110100101;
				8'b1001101: c <= 9'b100000100;
				8'b111111: c <= 9'b101000111;
				8'b1101110: c <= 9'b101000101;
				8'b1111011: c <= 9'b100111;
				8'b1001011: c <= 9'b111111000;
				8'b1101111: c <= 9'b11000010;
				8'b1101000: c <= 9'b1010011;
				8'b101100: c <= 9'b111100;
				8'b100100: c <= 9'b111010110;
				8'b1111000: c <= 9'b111100000;
				8'b1000101: c <= 9'b11110110;
				8'b1011001: c <= 9'b1011100;
				8'b110100: c <= 9'b11011111;
				8'b1111001: c <= 9'b111111111;
				8'b1110001: c <= 9'b1110100;
				8'b1001111: c <= 9'b110010100;
				8'b1100101: c <= 9'b110001111;
				8'b1111110: c <= 9'b110001010;
				8'b1111100: c <= 9'b11001010;
				8'b1010110: c <= 9'b111100011;
				8'b110010: c <= 9'b1001111;
				8'b1101101: c <= 9'b11100011;
				8'b100011: c <= 9'b1110010;
				8'b1110101: c <= 9'b10010110;
				8'b1111101: c <= 9'b11001;
				8'b101001: c <= 9'b111010000;
				8'b1010010: c <= 9'b110000000;
				8'b1011000: c <= 9'b110011011;
				8'b101110: c <= 9'b11000110;
				8'b1000001: c <= 9'b111111110;
				default: c <= 9'b0;
			endcase
			9'b11011111 : case(di)
				8'b1000011: c <= 9'b110011011;
				8'b101000: c <= 9'b111100010;
				8'b111010: c <= 9'b101101001;
				8'b110110: c <= 9'b110101001;
				8'b1100100: c <= 9'b110111000;
				8'b1000000: c <= 9'b111010110;
				8'b1110110: c <= 9'b11010010;
				8'b100101: c <= 9'b110010111;
				8'b101111: c <= 9'b110001110;
				8'b100110: c <= 9'b11111110;
				8'b1100011: c <= 9'b111110000;
				8'b1001000: c <= 9'b111000;
				8'b111000: c <= 9'b101101100;
				8'b110001: c <= 9'b101011011;
				8'b1010111: c <= 9'b110101110;
				8'b1001110: c <= 9'b111110000;
				8'b1101010: c <= 9'b11110011;
				8'b1001001: c <= 9'b111101000;
				8'b1100000: c <= 9'b101101101;
				8'b110111: c <= 9'b1110011;
				8'b1011101: c <= 9'b1001100;
				8'b1011011: c <= 9'b111110101;
				8'b111001: c <= 9'b101101100;
				8'b1001010: c <= 9'b111010110;
				8'b110011: c <= 9'b10010100;
				8'b1101100: c <= 9'b110111;
				8'b1110111: c <= 9'b100101100;
				8'b101011: c <= 9'b111110110;
				8'b1101011: c <= 9'b111010010;
				8'b111100: c <= 9'b1001100;
				8'b1000111: c <= 9'b100001010;
				8'b1011111: c <= 9'b10111010;
				8'b1110100: c <= 9'b110010000;
				8'b101101: c <= 9'b111001000;
				8'b1010011: c <= 9'b1110001;
				8'b1100001: c <= 9'b100101011;
				8'b110101: c <= 9'b111010100;
				8'b1000100: c <= 9'b111111011;
				8'b1010001: c <= 9'b101001;
				8'b1010100: c <= 9'b1010001;
				8'b1100110: c <= 9'b111001000;
				8'b101010: c <= 9'b111101110;
				8'b1011110: c <= 9'b11101101;
				8'b1100111: c <= 9'b100101111;
				8'b1011010: c <= 9'b11110111;
				8'b1000010: c <= 9'b10000111;
				8'b111101: c <= 9'b100110011;
				8'b110000: c <= 9'b111110000;
				8'b111110: c <= 9'b11001;
				8'b1100010: c <= 9'b100010000;
				8'b1110000: c <= 9'b11001010;
				8'b1101001: c <= 9'b10101000;
				8'b1110011: c <= 9'b111110110;
				8'b1001100: c <= 9'b111101010;
				8'b100001: c <= 9'b1011000;
				8'b1000110: c <= 9'b100011101;
				8'b1110010: c <= 9'b100110100;
				8'b1010000: c <= 9'b101010101;
				8'b1111010: c <= 9'b1001100;
				8'b1010101: c <= 9'b111100001;
				8'b111011: c <= 9'b110100010;
				8'b1001101: c <= 9'b100111101;
				8'b111111: c <= 9'b11;
				8'b1101110: c <= 9'b111001;
				8'b1111011: c <= 9'b110000111;
				8'b1001011: c <= 9'b1000;
				8'b1101111: c <= 9'b110000001;
				8'b1101000: c <= 9'b110001101;
				8'b101100: c <= 9'b10101;
				8'b100100: c <= 9'b11100110;
				8'b1111000: c <= 9'b101110;
				8'b1000101: c <= 9'b11101011;
				8'b1011001: c <= 9'b101101010;
				8'b110100: c <= 9'b110010011;
				8'b1111001: c <= 9'b101111010;
				8'b1110001: c <= 9'b100001;
				8'b1001111: c <= 9'b101001001;
				8'b1100101: c <= 9'b100110101;
				8'b1111110: c <= 9'b10100101;
				8'b1111100: c <= 9'b101000;
				8'b1010110: c <= 9'b10011001;
				8'b110010: c <= 9'b111000101;
				8'b1101101: c <= 9'b100111100;
				8'b100011: c <= 9'b1000101;
				8'b1110101: c <= 9'b10101100;
				8'b1111101: c <= 9'b10100011;
				8'b101001: c <= 9'b11001011;
				8'b1010010: c <= 9'b100110100;
				8'b1011000: c <= 9'b1010110;
				8'b101110: c <= 9'b111010111;
				8'b1000001: c <= 9'b111001010;
				default: c <= 9'b0;
			endcase
			9'b110010000 : case(di)
				8'b1000011: c <= 9'b1110111;
				8'b101000: c <= 9'b100100001;
				8'b111010: c <= 9'b101001001;
				8'b110110: c <= 9'b11110011;
				8'b1100100: c <= 9'b111110110;
				8'b1000000: c <= 9'b1000101;
				8'b1110110: c <= 9'b111111000;
				8'b100101: c <= 9'b10010000;
				8'b101111: c <= 9'b101001110;
				8'b100110: c <= 9'b10110101;
				8'b1100011: c <= 9'b101;
				8'b1001000: c <= 9'b101100101;
				8'b111000: c <= 9'b1100011;
				8'b110001: c <= 9'b111100111;
				8'b1010111: c <= 9'b10100;
				8'b1001110: c <= 9'b110001100;
				8'b1101010: c <= 9'b110011100;
				8'b1001001: c <= 9'b100100011;
				8'b1100000: c <= 9'b10110110;
				8'b110111: c <= 9'b11011000;
				8'b1011101: c <= 9'b1101110;
				8'b1011011: c <= 9'b10110111;
				8'b111001: c <= 9'b100010111;
				8'b1001010: c <= 9'b11011000;
				8'b110011: c <= 9'b111010001;
				8'b1101100: c <= 9'b10000110;
				8'b1110111: c <= 9'b1110100;
				8'b101011: c <= 9'b10111101;
				8'b1101011: c <= 9'b101110110;
				8'b111100: c <= 9'b10001011;
				8'b1000111: c <= 9'b1001001;
				8'b1011111: c <= 9'b110000;
				8'b1110100: c <= 9'b110111111;
				8'b101101: c <= 9'b10001011;
				8'b1010011: c <= 9'b1010000;
				8'b1100001: c <= 9'b101;
				8'b110101: c <= 9'b111000110;
				8'b1000100: c <= 9'b101101;
				8'b1010001: c <= 9'b1001011;
				8'b1010100: c <= 9'b11100101;
				8'b1100110: c <= 9'b100011001;
				8'b101010: c <= 9'b10101111;
				8'b1011110: c <= 9'b101010000;
				8'b1100111: c <= 9'b111000010;
				8'b1011010: c <= 9'b10101;
				8'b1000010: c <= 9'b110100011;
				8'b111101: c <= 9'b10100011;
				8'b110000: c <= 9'b1011101;
				8'b111110: c <= 9'b11010100;
				8'b1100010: c <= 9'b111111111;
				8'b1110000: c <= 9'b10111;
				8'b1101001: c <= 9'b111101101;
				8'b1110011: c <= 9'b100010110;
				8'b1001100: c <= 9'b110111111;
				8'b100001: c <= 9'b1111101;
				8'b1000110: c <= 9'b101011101;
				8'b1110010: c <= 9'b100;
				8'b1010000: c <= 9'b101111000;
				8'b1111010: c <= 9'b111100100;
				8'b1010101: c <= 9'b101100111;
				8'b111011: c <= 9'b110010001;
				8'b1001101: c <= 9'b101001110;
				8'b111111: c <= 9'b111111;
				8'b1101110: c <= 9'b110101;
				8'b1111011: c <= 9'b110001010;
				8'b1001011: c <= 9'b101110011;
				8'b1101111: c <= 9'b100000111;
				8'b1101000: c <= 9'b101001001;
				8'b101100: c <= 9'b10111010;
				8'b100100: c <= 9'b1011010;
				8'b1111000: c <= 9'b101111110;
				8'b1000101: c <= 9'b111000100;
				8'b1011001: c <= 9'b101010110;
				8'b110100: c <= 9'b11001010;
				8'b1111001: c <= 9'b10100100;
				8'b1110001: c <= 9'b10001011;
				8'b1001111: c <= 9'b111101111;
				8'b1100101: c <= 9'b11100011;
				8'b1111110: c <= 9'b110010101;
				8'b1111100: c <= 9'b11011101;
				8'b1010110: c <= 9'b111111;
				8'b110010: c <= 9'b100000110;
				8'b1101101: c <= 9'b111101;
				8'b100011: c <= 9'b1001010;
				8'b1110101: c <= 9'b110000010;
				8'b1111101: c <= 9'b100011111;
				8'b101001: c <= 9'b101001010;
				8'b1010010: c <= 9'b101011111;
				8'b1011000: c <= 9'b10101111;
				8'b101110: c <= 9'b110010111;
				8'b1000001: c <= 9'b10010;
				default: c <= 9'b0;
			endcase
			9'b1011101 : case(di)
				8'b1000011: c <= 9'b111000011;
				8'b101000: c <= 9'b110101010;
				8'b111010: c <= 9'b1110111;
				8'b110110: c <= 9'b10101110;
				8'b1100100: c <= 9'b10000111;
				8'b1000000: c <= 9'b110100100;
				8'b1110110: c <= 9'b11011001;
				8'b100101: c <= 9'b100011000;
				8'b101111: c <= 9'b111011001;
				8'b100110: c <= 9'b110011100;
				8'b1100011: c <= 9'b10010111;
				8'b1001000: c <= 9'b110110101;
				8'b111000: c <= 9'b100100110;
				8'b110001: c <= 9'b110000111;
				8'b1010111: c <= 9'b11101;
				8'b1001110: c <= 9'b11111;
				8'b1101010: c <= 9'b110110111;
				8'b1001001: c <= 9'b111100110;
				8'b1100000: c <= 9'b100000100;
				8'b110111: c <= 9'b111110101;
				8'b1011101: c <= 9'b11110001;
				8'b1011011: c <= 9'b1000100;
				8'b111001: c <= 9'b100001111;
				8'b1001010: c <= 9'b110100001;
				8'b110011: c <= 9'b101111010;
				8'b1101100: c <= 9'b111001001;
				8'b1110111: c <= 9'b110110010;
				8'b101011: c <= 9'b101010000;
				8'b1101011: c <= 9'b10011111;
				8'b111100: c <= 9'b10011101;
				8'b1000111: c <= 9'b11111001;
				8'b1011111: c <= 9'b110000010;
				8'b1110100: c <= 9'b1100000;
				8'b101101: c <= 9'b1101100;
				8'b1010011: c <= 9'b1100011;
				8'b1100001: c <= 9'b111100101;
				8'b110101: c <= 9'b110001000;
				8'b1000100: c <= 9'b10010001;
				8'b1010001: c <= 9'b11011;
				8'b1010100: c <= 9'b1011;
				8'b1100110: c <= 9'b11010;
				8'b101010: c <= 9'b101100011;
				8'b1011110: c <= 9'b101001011;
				8'b1100111: c <= 9'b1010010;
				8'b1011010: c <= 9'b100110011;
				8'b1000010: c <= 9'b100111010;
				8'b111101: c <= 9'b100010000;
				8'b110000: c <= 9'b100010110;
				8'b111110: c <= 9'b10011;
				8'b1100010: c <= 9'b1110101;
				8'b1110000: c <= 9'b110001101;
				8'b1101001: c <= 9'b110101110;
				8'b1110011: c <= 9'b110110000;
				8'b1001100: c <= 9'b110000101;
				8'b100001: c <= 9'b10111100;
				8'b1000110: c <= 9'b100010;
				8'b1110010: c <= 9'b11000101;
				8'b1010000: c <= 9'b1000;
				8'b1111010: c <= 9'b111001111;
				8'b1010101: c <= 9'b10011001;
				8'b111011: c <= 9'b101001000;
				8'b1001101: c <= 9'b101101010;
				8'b111111: c <= 9'b111011;
				8'b1101110: c <= 9'b110000000;
				8'b1111011: c <= 9'b110011101;
				8'b1001011: c <= 9'b10100111;
				8'b1101111: c <= 9'b101101001;
				8'b1101000: c <= 9'b1101101;
				8'b101100: c <= 9'b101101111;
				8'b100100: c <= 9'b1101111;
				8'b1111000: c <= 9'b1011001;
				8'b1000101: c <= 9'b100110011;
				8'b1011001: c <= 9'b101011110;
				8'b110100: c <= 9'b100100000;
				8'b1111001: c <= 9'b101011010;
				8'b1110001: c <= 9'b111001110;
				8'b1001111: c <= 9'b110101111;
				8'b1100101: c <= 9'b100101100;
				8'b1111110: c <= 9'b101100000;
				8'b1111100: c <= 9'b101010010;
				8'b1010110: c <= 9'b101110010;
				8'b110010: c <= 9'b111101101;
				8'b1101101: c <= 9'b10111000;
				8'b100011: c <= 9'b1001100;
				8'b1110101: c <= 9'b10111000;
				8'b1111101: c <= 9'b101101011;
				8'b101001: c <= 9'b10111100;
				8'b1010010: c <= 9'b1111011;
				8'b1011000: c <= 9'b101101001;
				8'b101110: c <= 9'b1110011;
				8'b1000001: c <= 9'b101110001;
				default: c <= 9'b0;
			endcase
			9'b11000101 : case(di)
				8'b1000011: c <= 9'b10110110;
				8'b101000: c <= 9'b11000111;
				8'b111010: c <= 9'b11110111;
				8'b110110: c <= 9'b100101111;
				8'b1100100: c <= 9'b110111100;
				8'b1000000: c <= 9'b1011;
				8'b1110110: c <= 9'b101110100;
				8'b100101: c <= 9'b10011001;
				8'b101111: c <= 9'b10100010;
				8'b100110: c <= 9'b1100100;
				8'b1100011: c <= 9'b11111100;
				8'b1001000: c <= 9'b111000111;
				8'b111000: c <= 9'b11000110;
				8'b110001: c <= 9'b11000011;
				8'b1010111: c <= 9'b1100111;
				8'b1001110: c <= 9'b10100011;
				8'b1101010: c <= 9'b110000111;
				8'b1001001: c <= 9'b1000010;
				8'b1100000: c <= 9'b11;
				8'b110111: c <= 9'b10001001;
				8'b1011101: c <= 9'b10;
				8'b1011011: c <= 9'b1100001;
				8'b111001: c <= 9'b110010100;
				8'b1001010: c <= 9'b11111100;
				8'b110011: c <= 9'b101001001;
				8'b1101100: c <= 9'b101101100;
				8'b1110111: c <= 9'b10110001;
				8'b101011: c <= 9'b111010100;
				8'b1101011: c <= 9'b110000000;
				8'b111100: c <= 9'b11111000;
				8'b1000111: c <= 9'b111000010;
				8'b1011111: c <= 9'b111111100;
				8'b1110100: c <= 9'b111111101;
				8'b101101: c <= 9'b100100011;
				8'b1010011: c <= 9'b1111101;
				8'b1100001: c <= 9'b101001000;
				8'b110101: c <= 9'b110101001;
				8'b1000100: c <= 9'b111111;
				8'b1010001: c <= 9'b1110100;
				8'b1010100: c <= 9'b110000010;
				8'b1100110: c <= 9'b110101110;
				8'b101010: c <= 9'b110111001;
				8'b1011110: c <= 9'b101100100;
				8'b1100111: c <= 9'b101001110;
				8'b1011010: c <= 9'b111100111;
				8'b1000010: c <= 9'b101100011;
				8'b111101: c <= 9'b1100001;
				8'b110000: c <= 9'b100101011;
				8'b111110: c <= 9'b1010110;
				8'b1100010: c <= 9'b101011000;
				8'b1110000: c <= 9'b1100000;
				8'b1101001: c <= 9'b11001010;
				8'b1110011: c <= 9'b10001011;
				8'b1001100: c <= 9'b110001;
				8'b100001: c <= 9'b1101111;
				8'b1000110: c <= 9'b100111001;
				8'b1110010: c <= 9'b100110101;
				8'b1010000: c <= 9'b111100010;
				8'b1111010: c <= 9'b11010;
				8'b1010101: c <= 9'b1;
				8'b111011: c <= 9'b100010111;
				8'b1001101: c <= 9'b111100011;
				8'b111111: c <= 9'b110100000;
				8'b1101110: c <= 9'b110110011;
				8'b1111011: c <= 9'b11001111;
				8'b1001011: c <= 9'b110101101;
				8'b1101111: c <= 9'b110;
				8'b1101000: c <= 9'b1111;
				8'b101100: c <= 9'b110101100;
				8'b100100: c <= 9'b10010000;
				8'b1111000: c <= 9'b11011001;
				8'b1000101: c <= 9'b100010111;
				8'b1011001: c <= 9'b110111100;
				8'b110100: c <= 9'b111011;
				8'b1111001: c <= 9'b101101000;
				8'b1110001: c <= 9'b1110101;
				8'b1001111: c <= 9'b101010010;
				8'b1100101: c <= 9'b110010100;
				8'b1111110: c <= 9'b1100000;
				8'b1111100: c <= 9'b110011110;
				8'b1010110: c <= 9'b111011001;
				8'b110010: c <= 9'b100111100;
				8'b1101101: c <= 9'b110100110;
				8'b100011: c <= 9'b11100000;
				8'b1110101: c <= 9'b11011110;
				8'b1111101: c <= 9'b110011101;
				8'b101001: c <= 9'b110111100;
				8'b1010010: c <= 9'b110000101;
				8'b1011000: c <= 9'b111010110;
				8'b101110: c <= 9'b101100110;
				8'b1000001: c <= 9'b110101011;
				default: c <= 9'b0;
			endcase
			9'b111111100 : case(di)
				8'b1000011: c <= 9'b100001011;
				8'b101000: c <= 9'b10110;
				8'b111010: c <= 9'b100011011;
				8'b110110: c <= 9'b11010000;
				8'b1100100: c <= 9'b1100;
				8'b1000000: c <= 9'b111010010;
				8'b1110110: c <= 9'b1110101;
				8'b100101: c <= 9'b11001101;
				8'b101111: c <= 9'b10101;
				8'b100110: c <= 9'b1010001;
				8'b1100011: c <= 9'b111010000;
				8'b1001000: c <= 9'b101101010;
				8'b111000: c <= 9'b100010101;
				8'b110001: c <= 9'b1111011;
				8'b1010111: c <= 9'b110;
				8'b1001110: c <= 9'b11101001;
				8'b1101010: c <= 9'b111001100;
				8'b1001001: c <= 9'b101100000;
				8'b1100000: c <= 9'b11110101;
				8'b110111: c <= 9'b100110111;
				8'b1011101: c <= 9'b101011111;
				8'b1011011: c <= 9'b110000111;
				8'b111001: c <= 9'b11010011;
				8'b1001010: c <= 9'b110010101;
				8'b110011: c <= 9'b1111000;
				8'b1101100: c <= 9'b101000010;
				8'b1110111: c <= 9'b11011010;
				8'b101011: c <= 9'b110101;
				8'b1101011: c <= 9'b10001101;
				8'b111100: c <= 9'b10101100;
				8'b1000111: c <= 9'b11000100;
				8'b1011111: c <= 9'b10100111;
				8'b1110100: c <= 9'b1000111;
				8'b101101: c <= 9'b11011010;
				8'b1010011: c <= 9'b110111000;
				8'b1100001: c <= 9'b110100;
				8'b110101: c <= 9'b11111100;
				8'b1000100: c <= 9'b11001110;
				8'b1010001: c <= 9'b100;
				8'b1010100: c <= 9'b10001110;
				8'b1100110: c <= 9'b1011111;
				8'b101010: c <= 9'b101110;
				8'b1011110: c <= 9'b10110100;
				8'b1100111: c <= 9'b101101010;
				8'b1011010: c <= 9'b111111110;
				8'b1000010: c <= 9'b1000;
				8'b111101: c <= 9'b1010010;
				8'b110000: c <= 9'b11111111;
				8'b111110: c <= 9'b100001001;
				8'b1100010: c <= 9'b111;
				8'b1110000: c <= 9'b111110001;
				8'b1101001: c <= 9'b10000111;
				8'b1110011: c <= 9'b111000100;
				8'b1001100: c <= 9'b11011001;
				8'b100001: c <= 9'b111000;
				8'b1000110: c <= 9'b111101001;
				8'b1110010: c <= 9'b101010010;
				8'b1010000: c <= 9'b11011101;
				8'b1111010: c <= 9'b100111;
				8'b1010101: c <= 9'b110100110;
				8'b111011: c <= 9'b111000010;
				8'b1001101: c <= 9'b111110001;
				8'b111111: c <= 9'b1011010;
				8'b1101110: c <= 9'b1001111;
				8'b1111011: c <= 9'b1100110;
				8'b1001011: c <= 9'b111111111;
				8'b1101111: c <= 9'b101110010;
				8'b1101000: c <= 9'b10111011;
				8'b101100: c <= 9'b101100111;
				8'b100100: c <= 9'b1010110;
				8'b1111000: c <= 9'b111101001;
				8'b1000101: c <= 9'b110010010;
				8'b1011001: c <= 9'b10001110;
				8'b110100: c <= 9'b101000110;
				8'b1111001: c <= 9'b10111111;
				8'b1110001: c <= 9'b110011010;
				8'b1001111: c <= 9'b10000000;
				8'b1100101: c <= 9'b10010111;
				8'b1111110: c <= 9'b11101000;
				8'b1111100: c <= 9'b10111110;
				8'b1010110: c <= 9'b11111110;
				8'b110010: c <= 9'b110111;
				8'b1101101: c <= 9'b111100100;
				8'b100011: c <= 9'b100110010;
				8'b1110101: c <= 9'b110111010;
				8'b1111101: c <= 9'b10001100;
				8'b101001: c <= 9'b101001001;
				8'b1010010: c <= 9'b1111100;
				8'b1011000: c <= 9'b1011011;
				8'b101110: c <= 9'b1011010;
				8'b1000001: c <= 9'b100010010;
				default: c <= 9'b0;
			endcase
			9'b11111111 : case(di)
				8'b1000011: c <= 9'b100101010;
				8'b101000: c <= 9'b11001;
				8'b111010: c <= 9'b11011;
				8'b110110: c <= 9'b1010111;
				8'b1100100: c <= 9'b111111101;
				8'b1000000: c <= 9'b101010011;
				8'b1110110: c <= 9'b111100010;
				8'b100101: c <= 9'b11001100;
				8'b101111: c <= 9'b111110001;
				8'b100110: c <= 9'b1100110;
				8'b1100011: c <= 9'b10110110;
				8'b1001000: c <= 9'b10101;
				8'b111000: c <= 9'b11001001;
				8'b110001: c <= 9'b10101100;
				8'b1010111: c <= 9'b10100100;
				8'b1001110: c <= 9'b110001;
				8'b1101010: c <= 9'b110111111;
				8'b1001001: c <= 9'b100010001;
				8'b1100000: c <= 9'b11110110;
				8'b110111: c <= 9'b101010011;
				8'b1011101: c <= 9'b110100110;
				8'b1011011: c <= 9'b111011100;
				8'b111001: c <= 9'b111011101;
				8'b1001010: c <= 9'b101111010;
				8'b110011: c <= 9'b11101111;
				8'b1101100: c <= 9'b10110011;
				8'b1110111: c <= 9'b1100000;
				8'b101011: c <= 9'b101011110;
				8'b1101011: c <= 9'b110;
				8'b111100: c <= 9'b111011100;
				8'b1000111: c <= 9'b110001000;
				8'b1011111: c <= 9'b111011;
				8'b1110100: c <= 9'b110000001;
				8'b101101: c <= 9'b1101000;
				8'b1010011: c <= 9'b100110100;
				8'b1100001: c <= 9'b100001011;
				8'b110101: c <= 9'b101001100;
				8'b1000100: c <= 9'b110111100;
				8'b1010001: c <= 9'b1100101;
				8'b1010100: c <= 9'b1000001;
				8'b1100110: c <= 9'b11000111;
				8'b101010: c <= 9'b100010;
				8'b1011110: c <= 9'b11011101;
				8'b1100111: c <= 9'b110011;
				8'b1011010: c <= 9'b110001100;
				8'b1000010: c <= 9'b10001101;
				8'b111101: c <= 9'b111001011;
				8'b110000: c <= 9'b100011000;
				8'b111110: c <= 9'b1000100;
				8'b1100010: c <= 9'b10011011;
				8'b1110000: c <= 9'b10100000;
				8'b1101001: c <= 9'b10110;
				8'b1110011: c <= 9'b11111010;
				8'b1001100: c <= 9'b1110010;
				8'b100001: c <= 9'b101100011;
				8'b1000110: c <= 9'b100100000;
				8'b1110010: c <= 9'b101111101;
				8'b1010000: c <= 9'b11000010;
				8'b1111010: c <= 9'b11111011;
				8'b1010101: c <= 9'b11110;
				8'b111011: c <= 9'b100101011;
				8'b1001101: c <= 9'b11100001;
				8'b111111: c <= 9'b100110111;
				8'b1101110: c <= 9'b100100000;
				8'b1111011: c <= 9'b101011;
				8'b1001011: c <= 9'b1010000;
				8'b1101111: c <= 9'b11111001;
				8'b1101000: c <= 9'b11000;
				8'b101100: c <= 9'b101001100;
				8'b100100: c <= 9'b100110;
				8'b1111000: c <= 9'b100100111;
				8'b1000101: c <= 9'b110111011;
				8'b1011001: c <= 9'b101001;
				8'b110100: c <= 9'b100010011;
				8'b1111001: c <= 9'b11011001;
				8'b1110001: c <= 9'b11111100;
				8'b1001111: c <= 9'b100101010;
				8'b1100101: c <= 9'b101001011;
				8'b1111110: c <= 9'b111100111;
				8'b1111100: c <= 9'b110011101;
				8'b1010110: c <= 9'b101100011;
				8'b110010: c <= 9'b11111000;
				8'b1101101: c <= 9'b111111;
				8'b100011: c <= 9'b1011110;
				8'b1110101: c <= 9'b1100100;
				8'b1111101: c <= 9'b111000010;
				8'b101001: c <= 9'b10111010;
				8'b1010010: c <= 9'b110101;
				8'b1011000: c <= 9'b111110011;
				8'b101110: c <= 9'b1011010;
				8'b1000001: c <= 9'b101000101;
				default: c <= 9'b0;
			endcase
			9'b101111101 : case(di)
				8'b1000011: c <= 9'b11010011;
				8'b101000: c <= 9'b101101000;
				8'b111010: c <= 9'b1001101;
				8'b110110: c <= 9'b100001101;
				8'b1100100: c <= 9'b1111;
				8'b1000000: c <= 9'b11011001;
				8'b1110110: c <= 9'b1100;
				8'b100101: c <= 9'b11100110;
				8'b101111: c <= 9'b11110110;
				8'b100110: c <= 9'b11011;
				8'b1100011: c <= 9'b111010110;
				8'b1001000: c <= 9'b11100100;
				8'b111000: c <= 9'b100010100;
				8'b110001: c <= 9'b111111000;
				8'b1010111: c <= 9'b110100110;
				8'b1001110: c <= 9'b11110100;
				8'b1101010: c <= 9'b100111110;
				8'b1001001: c <= 9'b111100001;
				8'b1100000: c <= 9'b10100000;
				8'b110111: c <= 9'b11111;
				8'b1011101: c <= 9'b100110110;
				8'b1011011: c <= 9'b1011000;
				8'b111001: c <= 9'b101100000;
				8'b1001010: c <= 9'b111111110;
				8'b110011: c <= 9'b110011;
				8'b1101100: c <= 9'b111000;
				8'b1110111: c <= 9'b1010111;
				8'b101011: c <= 9'b100000011;
				8'b1101011: c <= 9'b100110000;
				8'b111100: c <= 9'b1000111;
				8'b1000111: c <= 9'b101101101;
				8'b1011111: c <= 9'b111010101;
				8'b1110100: c <= 9'b110111010;
				8'b101101: c <= 9'b100111011;
				8'b1010011: c <= 9'b10001000;
				8'b1100001: c <= 9'b111000100;
				8'b110101: c <= 9'b100011101;
				8'b1000100: c <= 9'b110001010;
				8'b1010001: c <= 9'b101000110;
				8'b1010100: c <= 9'b111011011;
				8'b1100110: c <= 9'b110;
				8'b101010: c <= 9'b100011011;
				8'b1011110: c <= 9'b101000101;
				8'b1100111: c <= 9'b10110;
				8'b1011010: c <= 9'b101010001;
				8'b1000010: c <= 9'b101000101;
				8'b111101: c <= 9'b111011011;
				8'b110000: c <= 9'b10100011;
				8'b111110: c <= 9'b11111001;
				8'b1100010: c <= 9'b100100011;
				8'b1110000: c <= 9'b11010100;
				8'b1101001: c <= 9'b11001010;
				8'b1110011: c <= 9'b11011010;
				8'b1001100: c <= 9'b101110011;
				8'b100001: c <= 9'b11000100;
				8'b1000110: c <= 9'b10001101;
				8'b1110010: c <= 9'b100000101;
				8'b1010000: c <= 9'b10111001;
				8'b1111010: c <= 9'b1000001;
				8'b1010101: c <= 9'b110000001;
				8'b111011: c <= 9'b100100111;
				8'b1001101: c <= 9'b11110101;
				8'b111111: c <= 9'b101000010;
				8'b1101110: c <= 9'b1100011;
				8'b1111011: c <= 9'b100110011;
				8'b1001011: c <= 9'b111110011;
				8'b1101111: c <= 9'b100001011;
				8'b1101000: c <= 9'b1111100;
				8'b101100: c <= 9'b101001100;
				8'b100100: c <= 9'b110010;
				8'b1111000: c <= 9'b10110110;
				8'b1000101: c <= 9'b110011101;
				8'b1011001: c <= 9'b111110000;
				8'b110100: c <= 9'b111111011;
				8'b1111001: c <= 9'b101011110;
				8'b1110001: c <= 9'b100100101;
				8'b1001111: c <= 9'b111011101;
				8'b1100101: c <= 9'b110110011;
				8'b1111110: c <= 9'b110110111;
				8'b1111100: c <= 9'b110000110;
				8'b1010110: c <= 9'b1011010;
				8'b110010: c <= 9'b101111110;
				8'b1101101: c <= 9'b100000111;
				8'b100011: c <= 9'b111001110;
				8'b1110101: c <= 9'b11110010;
				8'b1111101: c <= 9'b111011100;
				8'b101001: c <= 9'b10001010;
				8'b1010010: c <= 9'b111100000;
				8'b1011000: c <= 9'b10000011;
				8'b101110: c <= 9'b110111011;
				8'b1000001: c <= 9'b10111101;
				default: c <= 9'b0;
			endcase
			9'b111010101 : case(di)
				8'b1000011: c <= 9'b1011000;
				8'b101000: c <= 9'b101101100;
				8'b111010: c <= 9'b100001001;
				8'b110110: c <= 9'b100010010;
				8'b1100100: c <= 9'b100100011;
				8'b1000000: c <= 9'b10101011;
				8'b1110110: c <= 9'b100011000;
				8'b100101: c <= 9'b111111001;
				8'b101111: c <= 9'b101000111;
				8'b100110: c <= 9'b111011010;
				8'b1100011: c <= 9'b101110000;
				8'b1001000: c <= 9'b11110010;
				8'b111000: c <= 9'b1100011;
				8'b110001: c <= 9'b10101010;
				8'b1010111: c <= 9'b1;
				8'b1001110: c <= 9'b100100101;
				8'b1101010: c <= 9'b10111011;
				8'b1001001: c <= 9'b100111011;
				8'b1100000: c <= 9'b101010000;
				8'b110111: c <= 9'b100011010;
				8'b1011101: c <= 9'b110001101;
				8'b1011011: c <= 9'b110011101;
				8'b111001: c <= 9'b10000000;
				8'b1001010: c <= 9'b111101000;
				8'b110011: c <= 9'b10101011;
				8'b1101100: c <= 9'b110100;
				8'b1110111: c <= 9'b11100010;
				8'b101011: c <= 9'b100111011;
				8'b1101011: c <= 9'b101011001;
				8'b111100: c <= 9'b100110011;
				8'b1000111: c <= 9'b10100010;
				8'b1011111: c <= 9'b101100;
				8'b1110100: c <= 9'b100000011;
				8'b101101: c <= 9'b100101110;
				8'b1010011: c <= 9'b100000110;
				8'b1100001: c <= 9'b110101100;
				8'b110101: c <= 9'b11010010;
				8'b1000100: c <= 9'b101010000;
				8'b1010001: c <= 9'b11100011;
				8'b1010100: c <= 9'b10011011;
				8'b1100110: c <= 9'b111001000;
				8'b101010: c <= 9'b101100110;
				8'b1011110: c <= 9'b10101011;
				8'b1100111: c <= 9'b1011100;
				8'b1011010: c <= 9'b110010010;
				8'b1000010: c <= 9'b101110011;
				8'b111101: c <= 9'b11110011;
				8'b110000: c <= 9'b111001010;
				8'b111110: c <= 9'b10101110;
				8'b1100010: c <= 9'b1101001;
				8'b1110000: c <= 9'b101100111;
				8'b1101001: c <= 9'b1001110;
				8'b1110011: c <= 9'b101111;
				8'b1001100: c <= 9'b110100101;
				8'b100001: c <= 9'b10101;
				8'b1000110: c <= 9'b111000111;
				8'b1110010: c <= 9'b111000110;
				8'b1010000: c <= 9'b1110100;
				8'b1111010: c <= 9'b110000001;
				8'b1010101: c <= 9'b100010101;
				8'b111011: c <= 9'b11100;
				8'b1001101: c <= 9'b101001011;
				8'b111111: c <= 9'b100000100;
				8'b1101110: c <= 9'b111100110;
				8'b1111011: c <= 9'b100010;
				8'b1001011: c <= 9'b111101110;
				8'b1101111: c <= 9'b111101010;
				8'b1101000: c <= 9'b110000101;
				8'b101100: c <= 9'b100010;
				8'b100100: c <= 9'b110000111;
				8'b1111000: c <= 9'b110100110;
				8'b1000101: c <= 9'b101110010;
				8'b1011001: c <= 9'b110001010;
				8'b110100: c <= 9'b11001000;
				8'b1111001: c <= 9'b110010;
				8'b1110001: c <= 9'b111100111;
				8'b1001111: c <= 9'b111100110;
				8'b1100101: c <= 9'b111101000;
				8'b1111110: c <= 9'b111001000;
				8'b1111100: c <= 9'b10101110;
				8'b1010110: c <= 9'b1010001;
				8'b110010: c <= 9'b11111100;
				8'b1101101: c <= 9'b10000110;
				8'b100011: c <= 9'b111001011;
				8'b1110101: c <= 9'b1100011;
				8'b1111101: c <= 9'b11111011;
				8'b101001: c <= 9'b11001;
				8'b1010010: c <= 9'b110100001;
				8'b1011000: c <= 9'b11011100;
				8'b101110: c <= 9'b11001010;
				8'b1000001: c <= 9'b11010111;
				default: c <= 9'b0;
			endcase
			9'b101111 : case(di)
				8'b1000011: c <= 9'b111110011;
				8'b101000: c <= 9'b1010101;
				8'b111010: c <= 9'b101001;
				8'b110110: c <= 9'b1100001;
				8'b1100100: c <= 9'b10010111;
				8'b1000000: c <= 9'b11111000;
				8'b1110110: c <= 9'b11100000;
				8'b100101: c <= 9'b100010011;
				8'b101111: c <= 9'b10111101;
				8'b100110: c <= 9'b1101101;
				8'b1100011: c <= 9'b11100011;
				8'b1001000: c <= 9'b11010;
				8'b111000: c <= 9'b100011010;
				8'b110001: c <= 9'b100011001;
				8'b1010111: c <= 9'b1110011;
				8'b1001110: c <= 9'b10101111;
				8'b1101010: c <= 9'b111011;
				8'b1001001: c <= 9'b11010010;
				8'b1100000: c <= 9'b1111001;
				8'b110111: c <= 9'b10010101;
				8'b1011101: c <= 9'b100101100;
				8'b1011011: c <= 9'b110110000;
				8'b111001: c <= 9'b110101010;
				8'b1001010: c <= 9'b11100011;
				8'b110011: c <= 9'b10100111;
				8'b1101100: c <= 9'b11;
				8'b1110111: c <= 9'b101111110;
				8'b101011: c <= 9'b11010111;
				8'b1101011: c <= 9'b110011;
				8'b111100: c <= 9'b1100;
				8'b1000111: c <= 9'b110110010;
				8'b1011111: c <= 9'b11010011;
				8'b1110100: c <= 9'b111110100;
				8'b101101: c <= 9'b101100011;
				8'b1010011: c <= 9'b110001111;
				8'b1100001: c <= 9'b100011000;
				8'b110101: c <= 9'b100101110;
				8'b1000100: c <= 9'b100110000;
				8'b1010001: c <= 9'b11101011;
				8'b1010100: c <= 9'b1101111;
				8'b1100110: c <= 9'b1101100;
				8'b101010: c <= 9'b110001001;
				8'b1011110: c <= 9'b11010000;
				8'b1100111: c <= 9'b101010010;
				8'b1011010: c <= 9'b101110001;
				8'b1000010: c <= 9'b11110100;
				8'b111101: c <= 9'b11001000;
				8'b110000: c <= 9'b110111001;
				8'b111110: c <= 9'b10110;
				8'b1100010: c <= 9'b101010001;
				8'b1110000: c <= 9'b100110110;
				8'b1101001: c <= 9'b1011010;
				8'b1110011: c <= 9'b110100110;
				8'b1001100: c <= 9'b100001111;
				8'b100001: c <= 9'b11101111;
				8'b1000110: c <= 9'b110101100;
				8'b1110010: c <= 9'b11000;
				8'b1010000: c <= 9'b10011000;
				8'b1111010: c <= 9'b1110011;
				8'b1010101: c <= 9'b1010000;
				8'b111011: c <= 9'b110111110;
				8'b1001101: c <= 9'b100110110;
				8'b111111: c <= 9'b101001100;
				8'b1101110: c <= 9'b100110;
				8'b1111011: c <= 9'b101110001;
				8'b1001011: c <= 9'b1100001;
				8'b1101111: c <= 9'b111101110;
				8'b1101000: c <= 9'b10011101;
				8'b101100: c <= 9'b100010011;
				8'b100100: c <= 9'b101101000;
				8'b1111000: c <= 9'b101001110;
				8'b1000101: c <= 9'b10101010;
				8'b1011001: c <= 9'b110011101;
				8'b110100: c <= 9'b111010010;
				8'b1111001: c <= 9'b101010;
				8'b1110001: c <= 9'b111101101;
				8'b1001111: c <= 9'b10111101;
				8'b1100101: c <= 9'b110100000;
				8'b1111110: c <= 9'b101100010;
				8'b1111100: c <= 9'b101111010;
				8'b1010110: c <= 9'b110010011;
				8'b110010: c <= 9'b10100010;
				8'b1101101: c <= 9'b10011011;
				8'b100011: c <= 9'b110010011;
				8'b1110101: c <= 9'b10111011;
				8'b1111101: c <= 9'b11111010;
				8'b101001: c <= 9'b1101000;
				8'b1010010: c <= 9'b110000101;
				8'b1011000: c <= 9'b101111010;
				8'b101110: c <= 9'b10011011;
				8'b1000001: c <= 9'b100100000;
				default: c <= 9'b0;
			endcase
			9'b111110100 : case(di)
				8'b1000011: c <= 9'b1000;
				8'b101000: c <= 9'b110111001;
				8'b111010: c <= 9'b111011111;
				8'b110110: c <= 9'b100101000;
				8'b1100100: c <= 9'b10111100;
				8'b1000000: c <= 9'b11110110;
				8'b1110110: c <= 9'b11001;
				8'b100101: c <= 9'b111011111;
				8'b101111: c <= 9'b110111110;
				8'b100110: c <= 9'b110100011;
				8'b1100011: c <= 9'b100000100;
				8'b1001000: c <= 9'b11000111;
				8'b111000: c <= 9'b10100010;
				8'b110001: c <= 9'b11001011;
				8'b1010111: c <= 9'b11011100;
				8'b1001110: c <= 9'b1010111;
				8'b1101010: c <= 9'b100101001;
				8'b1001001: c <= 9'b101100010;
				8'b1100000: c <= 9'b1111;
				8'b110111: c <= 9'b110000010;
				8'b1011101: c <= 9'b110110;
				8'b1011011: c <= 9'b10010011;
				8'b111001: c <= 9'b1111;
				8'b1001010: c <= 9'b1001010;
				8'b110011: c <= 9'b101001111;
				8'b1101100: c <= 9'b10100000;
				8'b1110111: c <= 9'b11111110;
				8'b101011: c <= 9'b11101;
				8'b1101011: c <= 9'b1011;
				8'b111100: c <= 9'b110000110;
				8'b1000111: c <= 9'b10110011;
				8'b1011111: c <= 9'b100111000;
				8'b1110100: c <= 9'b1100010;
				8'b101101: c <= 9'b10100011;
				8'b1010011: c <= 9'b1101100;
				8'b1100001: c <= 9'b11011010;
				8'b110101: c <= 9'b100010011;
				8'b1000100: c <= 9'b1011001;
				8'b1010001: c <= 9'b110111100;
				8'b1010100: c <= 9'b111010010;
				8'b1100110: c <= 9'b101011000;
				8'b101010: c <= 9'b11001110;
				8'b1011110: c <= 9'b10011;
				8'b1100111: c <= 9'b110010101;
				8'b1011010: c <= 9'b110100110;
				8'b1000010: c <= 9'b1011010;
				8'b111101: c <= 9'b1110001;
				8'b110000: c <= 9'b101011011;
				8'b111110: c <= 9'b10110111;
				8'b1100010: c <= 9'b100000010;
				8'b1110000: c <= 9'b110011010;
				8'b1101001: c <= 9'b11111000;
				8'b1110011: c <= 9'b11010;
				8'b1001100: c <= 9'b111010001;
				8'b100001: c <= 9'b11110000;
				8'b1000110: c <= 9'b1011;
				8'b1110010: c <= 9'b11100010;
				8'b1010000: c <= 9'b11111;
				8'b1111010: c <= 9'b1010011;
				8'b1010101: c <= 9'b111000110;
				8'b111011: c <= 9'b10000101;
				8'b1001101: c <= 9'b1000010;
				8'b111111: c <= 9'b1010011;
				8'b1101110: c <= 9'b11101101;
				8'b1111011: c <= 9'b1100001;
				8'b1001011: c <= 9'b101000011;
				8'b1101111: c <= 9'b10100110;
				8'b1101000: c <= 9'b100100100;
				8'b101100: c <= 9'b10010000;
				8'b100100: c <= 9'b111;
				8'b1111000: c <= 9'b110000011;
				8'b1000101: c <= 9'b10011000;
				8'b1011001: c <= 9'b100011111;
				8'b110100: c <= 9'b100111100;
				8'b1111001: c <= 9'b111101100;
				8'b1110001: c <= 9'b101110011;
				8'b1001111: c <= 9'b111011111;
				8'b1100101: c <= 9'b1101010;
				8'b1111110: c <= 9'b11100101;
				8'b1111100: c <= 9'b111110001;
				8'b1010110: c <= 9'b101011010;
				8'b110010: c <= 9'b100000000;
				8'b1101101: c <= 9'b11001100;
				8'b100011: c <= 9'b100011111;
				8'b1110101: c <= 9'b110111001;
				8'b1111101: c <= 9'b11001100;
				8'b101001: c <= 9'b10100101;
				8'b1010010: c <= 9'b101001011;
				8'b1011000: c <= 9'b100001100;
				8'b101110: c <= 9'b1011100;
				8'b1000001: c <= 9'b11110001;
				default: c <= 9'b0;
			endcase
			9'b100100100 : case(di)
				8'b1000011: c <= 9'b101100101;
				8'b101000: c <= 9'b110100110;
				8'b111010: c <= 9'b11001111;
				8'b110110: c <= 9'b101011111;
				8'b1100100: c <= 9'b10001000;
				8'b1000000: c <= 9'b1011110;
				8'b1110110: c <= 9'b11011110;
				8'b100101: c <= 9'b11011101;
				8'b101111: c <= 9'b101100011;
				8'b100110: c <= 9'b10010001;
				8'b1100011: c <= 9'b110001;
				8'b1001000: c <= 9'b110101110;
				8'b111000: c <= 9'b101101111;
				8'b110001: c <= 9'b1100011;
				8'b1010111: c <= 9'b101011010;
				8'b1001110: c <= 9'b111101;
				8'b1101010: c <= 9'b110101100;
				8'b1001001: c <= 9'b10110011;
				8'b1100000: c <= 9'b11100000;
				8'b110111: c <= 9'b101000010;
				8'b1011101: c <= 9'b111011010;
				8'b1011011: c <= 9'b10010111;
				8'b111001: c <= 9'b101101;
				8'b1001010: c <= 9'b1110100;
				8'b110011: c <= 9'b110101101;
				8'b1101100: c <= 9'b10;
				8'b1110111: c <= 9'b110100;
				8'b101011: c <= 9'b111110101;
				8'b1101011: c <= 9'b110111011;
				8'b111100: c <= 9'b111010010;
				8'b1000111: c <= 9'b101100000;
				8'b1011111: c <= 9'b110010011;
				8'b1110100: c <= 9'b101101010;
				8'b101101: c <= 9'b10001010;
				8'b1010011: c <= 9'b111001010;
				8'b1100001: c <= 9'b111100000;
				8'b110101: c <= 9'b100100010;
				8'b1000100: c <= 9'b101101111;
				8'b1010001: c <= 9'b10111110;
				8'b1010100: c <= 9'b111;
				8'b1100110: c <= 9'b111010000;
				8'b101010: c <= 9'b1110011;
				8'b1011110: c <= 9'b10111100;
				8'b1100111: c <= 9'b100100;
				8'b1011010: c <= 9'b101110100;
				8'b1000010: c <= 9'b11111110;
				8'b111101: c <= 9'b100011010;
				8'b110000: c <= 9'b11010100;
				8'b111110: c <= 9'b11010100;
				8'b1100010: c <= 9'b1100100;
				8'b1110000: c <= 9'b11110;
				8'b1101001: c <= 9'b10000;
				8'b1110011: c <= 9'b11011001;
				8'b1001100: c <= 9'b1110001;
				8'b100001: c <= 9'b11000010;
				8'b1000110: c <= 9'b110010110;
				8'b1110010: c <= 9'b1101000;
				8'b1010000: c <= 9'b11100000;
				8'b1111010: c <= 9'b101001111;
				8'b1010101: c <= 9'b10111010;
				8'b111011: c <= 9'b101001010;
				8'b1001101: c <= 9'b11110010;
				8'b111111: c <= 9'b1101;
				8'b1101110: c <= 9'b100110110;
				8'b1111011: c <= 9'b10100111;
				8'b1001011: c <= 9'b11110001;
				8'b1101111: c <= 9'b1010101;
				8'b1101000: c <= 9'b100100110;
				8'b101100: c <= 9'b100010110;
				8'b100100: c <= 9'b111011010;
				8'b1111000: c <= 9'b10000000;
				8'b1000101: c <= 9'b110010110;
				8'b1011001: c <= 9'b110100000;
				8'b110100: c <= 9'b101101010;
				8'b1111001: c <= 9'b10100110;
				8'b1110001: c <= 9'b1110011;
				8'b1001111: c <= 9'b11001110;
				8'b1100101: c <= 9'b11111001;
				8'b1111110: c <= 9'b11101;
				8'b1111100: c <= 9'b100001;
				8'b1010110: c <= 9'b110011001;
				8'b110010: c <= 9'b111111010;
				8'b1101101: c <= 9'b100110000;
				8'b100011: c <= 9'b100101101;
				8'b1110101: c <= 9'b100111011;
				8'b1111101: c <= 9'b11010010;
				8'b101001: c <= 9'b1011;
				8'b1010010: c <= 9'b10010000;
				8'b1011000: c <= 9'b101001001;
				8'b101110: c <= 9'b1110110;
				8'b1000001: c <= 9'b110011111;
				default: c <= 9'b0;
			endcase
			9'b1110110 : case(di)
				8'b1000011: c <= 9'b101000;
				8'b101000: c <= 9'b1110000;
				8'b111010: c <= 9'b1110000;
				8'b110110: c <= 9'b1101101;
				8'b1100100: c <= 9'b101001100;
				8'b1000000: c <= 9'b110100001;
				8'b1110110: c <= 9'b111101111;
				8'b100101: c <= 9'b1010000;
				8'b101111: c <= 9'b111010110;
				8'b100110: c <= 9'b100110100;
				8'b1100011: c <= 9'b11010;
				8'b1001000: c <= 9'b110101101;
				8'b111000: c <= 9'b101010111;
				8'b110001: c <= 9'b11101000;
				8'b1010111: c <= 9'b111010010;
				8'b1001110: c <= 9'b1100110;
				8'b1101010: c <= 9'b110100011;
				8'b1001001: c <= 9'b11110111;
				8'b1100000: c <= 9'b10011001;
				8'b110111: c <= 9'b100001010;
				8'b1011101: c <= 9'b101010010;
				8'b1011011: c <= 9'b111101100;
				8'b111001: c <= 9'b1000001;
				8'b1001010: c <= 9'b110011101;
				8'b110011: c <= 9'b10010000;
				8'b1101100: c <= 9'b1100011;
				8'b1110111: c <= 9'b111111001;
				8'b101011: c <= 9'b10001011;
				8'b1101011: c <= 9'b1011111;
				8'b111100: c <= 9'b100011100;
				8'b1000111: c <= 9'b10110010;
				8'b1011111: c <= 9'b101010010;
				8'b1110100: c <= 9'b111110000;
				8'b101101: c <= 9'b10100101;
				8'b1010011: c <= 9'b111000;
				8'b1100001: c <= 9'b111011011;
				8'b110101: c <= 9'b100001100;
				8'b1000100: c <= 9'b11111011;
				8'b1010001: c <= 9'b110001000;
				8'b1010100: c <= 9'b110111111;
				8'b1100110: c <= 9'b101001001;
				8'b101010: c <= 9'b1101101;
				8'b1011110: c <= 9'b100100;
				8'b1100111: c <= 9'b1011010;
				8'b1011010: c <= 9'b101010011;
				8'b1000010: c <= 9'b111000100;
				8'b111101: c <= 9'b10011001;
				8'b110000: c <= 9'b100000000;
				8'b111110: c <= 9'b100110000;
				8'b1100010: c <= 9'b110100111;
				8'b1110000: c <= 9'b111011110;
				8'b1101001: c <= 9'b100000101;
				8'b1110011: c <= 9'b11001011;
				8'b1001100: c <= 9'b10110110;
				8'b100001: c <= 9'b110100011;
				8'b1000110: c <= 9'b100111000;
				8'b1110010: c <= 9'b1011100;
				8'b1010000: c <= 9'b11111110;
				8'b1111010: c <= 9'b111010100;
				8'b1010101: c <= 9'b1010010;
				8'b111011: c <= 9'b100010;
				8'b1001101: c <= 9'b101010;
				8'b111111: c <= 9'b10010100;
				8'b1101110: c <= 9'b101110100;
				8'b1111011: c <= 9'b11110011;
				8'b1001011: c <= 9'b1001111;
				8'b1101111: c <= 9'b11001000;
				8'b1101000: c <= 9'b111011001;
				8'b101100: c <= 9'b1001101;
				8'b100100: c <= 9'b111111101;
				8'b1111000: c <= 9'b100110000;
				8'b1000101: c <= 9'b11110010;
				8'b1011001: c <= 9'b11011001;
				8'b110100: c <= 9'b10111111;
				8'b1111001: c <= 9'b100111011;
				8'b1110001: c <= 9'b11011011;
				8'b1001111: c <= 9'b110010;
				8'b1100101: c <= 9'b11101101;
				8'b1111110: c <= 9'b10011101;
				8'b1111100: c <= 9'b101000110;
				8'b1010110: c <= 9'b1100100;
				8'b110010: c <= 9'b10000010;
				8'b1101101: c <= 9'b1011;
				8'b100011: c <= 9'b11010010;
				8'b1110101: c <= 9'b100101110;
				8'b1111101: c <= 9'b101111110;
				8'b101001: c <= 9'b10111011;
				8'b1010010: c <= 9'b100000000;
				8'b1011000: c <= 9'b1100010;
				8'b101110: c <= 9'b111010011;
				8'b1000001: c <= 9'b111100111;
				default: c <= 9'b0;
			endcase
			9'b111010011 : case(di)
				8'b1000011: c <= 9'b111111101;
				8'b101000: c <= 9'b11100111;
				8'b111010: c <= 9'b10111010;
				8'b110110: c <= 9'b111101110;
				8'b1100100: c <= 9'b1101101;
				8'b1000000: c <= 9'b111011;
				8'b1110110: c <= 9'b10100011;
				8'b100101: c <= 9'b100000100;
				8'b101111: c <= 9'b101001001;
				8'b100110: c <= 9'b101001;
				8'b1100011: c <= 9'b10011000;
				8'b1001000: c <= 9'b110010010;
				8'b111000: c <= 9'b101100110;
				8'b110001: c <= 9'b101100111;
				8'b1010111: c <= 9'b110010011;
				8'b1001110: c <= 9'b10010000;
				8'b1101010: c <= 9'b11111000;
				8'b1001001: c <= 9'b111100001;
				8'b1100000: c <= 9'b100010101;
				8'b110111: c <= 9'b100110110;
				8'b1011101: c <= 9'b1;
				8'b1011011: c <= 9'b110100100;
				8'b111001: c <= 9'b101010110;
				8'b1001010: c <= 9'b11011;
				8'b110011: c <= 9'b1010011;
				8'b1101100: c <= 9'b110011001;
				8'b1110111: c <= 9'b10100111;
				8'b101011: c <= 9'b11101;
				8'b1101011: c <= 9'b110111110;
				8'b111100: c <= 9'b1;
				8'b1000111: c <= 9'b11100100;
				8'b1011111: c <= 9'b111000000;
				8'b1110100: c <= 9'b10011100;
				8'b101101: c <= 9'b110011100;
				8'b1010011: c <= 9'b11010010;
				8'b1100001: c <= 9'b100100101;
				8'b110101: c <= 9'b11100110;
				8'b1000100: c <= 9'b111001110;
				8'b1010001: c <= 9'b1110;
				8'b1010100: c <= 9'b100110000;
				8'b1100110: c <= 9'b101000100;
				8'b101010: c <= 9'b10110010;
				8'b1011110: c <= 9'b1001110;
				8'b1100111: c <= 9'b111000;
				8'b1011010: c <= 9'b101001011;
				8'b1000010: c <= 9'b111010000;
				8'b111101: c <= 9'b101101;
				8'b110000: c <= 9'b111010110;
				8'b111110: c <= 9'b1000101;
				8'b1100010: c <= 9'b1000;
				8'b1110000: c <= 9'b110000111;
				8'b1101001: c <= 9'b111001001;
				8'b1110011: c <= 9'b110110010;
				8'b1001100: c <= 9'b10010001;
				8'b100001: c <= 9'b10000001;
				8'b1000110: c <= 9'b101101100;
				8'b1110010: c <= 9'b111010110;
				8'b1010000: c <= 9'b11100110;
				8'b1111010: c <= 9'b10101;
				8'b1010101: c <= 9'b101000;
				8'b111011: c <= 9'b100011001;
				8'b1001101: c <= 9'b100111000;
				8'b111111: c <= 9'b110000000;
				8'b1101110: c <= 9'b111100100;
				8'b1111011: c <= 9'b101010000;
				8'b1001011: c <= 9'b11010000;
				8'b1101111: c <= 9'b11101001;
				8'b1101000: c <= 9'b1110000;
				8'b101100: c <= 9'b100110100;
				8'b100100: c <= 9'b110110;
				8'b1111000: c <= 9'b110001001;
				8'b1000101: c <= 9'b100000100;
				8'b1011001: c <= 9'b100000111;
				8'b110100: c <= 9'b110101101;
				8'b1111001: c <= 9'b101010111;
				8'b1110001: c <= 9'b1000011;
				8'b1001111: c <= 9'b10000110;
				8'b1100101: c <= 9'b111111110;
				8'b1111110: c <= 9'b10011001;
				8'b1111100: c <= 9'b11011110;
				8'b1010110: c <= 9'b100011111;
				8'b110010: c <= 9'b101000100;
				8'b1101101: c <= 9'b10001110;
				8'b100011: c <= 9'b101001010;
				8'b1110101: c <= 9'b111010;
				8'b1111101: c <= 9'b11011101;
				8'b101001: c <= 9'b101111000;
				8'b1010010: c <= 9'b111011100;
				8'b1011000: c <= 9'b111111011;
				8'b101110: c <= 9'b101011100;
				8'b1000001: c <= 9'b110000011;
				default: c <= 9'b0;
			endcase
			9'b101011100 : case(di)
				8'b1000011: c <= 9'b11101100;
				8'b101000: c <= 9'b10001111;
				8'b111010: c <= 9'b110001110;
				8'b110110: c <= 9'b111010100;
				8'b1100100: c <= 9'b1110101;
				8'b1000000: c <= 9'b1110001;
				8'b1110110: c <= 9'b111100010;
				8'b100101: c <= 9'b111000101;
				8'b101111: c <= 9'b111100010;
				8'b100110: c <= 9'b11011;
				8'b1100011: c <= 9'b11111;
				8'b1001000: c <= 9'b11111010;
				8'b111000: c <= 9'b11001110;
				8'b110001: c <= 9'b110011000;
				8'b1010111: c <= 9'b1011000;
				8'b1001110: c <= 9'b11000011;
				8'b1101010: c <= 9'b10000111;
				8'b1001001: c <= 9'b1101001;
				8'b1100000: c <= 9'b110110011;
				8'b110111: c <= 9'b111100010;
				8'b1011101: c <= 9'b111000011;
				8'b1011011: c <= 9'b101000100;
				8'b111001: c <= 9'b10001100;
				8'b1001010: c <= 9'b110101110;
				8'b110011: c <= 9'b100110100;
				8'b1101100: c <= 9'b100110;
				8'b1110111: c <= 9'b1001011;
				8'b101011: c <= 9'b101101;
				8'b1101011: c <= 9'b100010011;
				8'b111100: c <= 9'b110101;
				8'b1000111: c <= 9'b10110011;
				8'b1011111: c <= 9'b10110010;
				8'b1110100: c <= 9'b1000010;
				8'b101101: c <= 9'b101001100;
				8'b1010011: c <= 9'b11111000;
				8'b1100001: c <= 9'b10110;
				8'b110101: c <= 9'b10100010;
				8'b1000100: c <= 9'b1010110;
				8'b1010001: c <= 9'b11010;
				8'b1010100: c <= 9'b1001010;
				8'b1100110: c <= 9'b1001110;
				8'b101010: c <= 9'b1101101;
				8'b1011110: c <= 9'b10100000;
				8'b1100111: c <= 9'b111101111;
				8'b1011010: c <= 9'b110010110;
				8'b1000010: c <= 9'b10010001;
				8'b111101: c <= 9'b110000111;
				8'b110000: c <= 9'b10100111;
				8'b111110: c <= 9'b1000010;
				8'b1100010: c <= 9'b111100010;
				8'b1110000: c <= 9'b1011010;
				8'b1101001: c <= 9'b100101111;
				8'b1110011: c <= 9'b110101010;
				8'b1001100: c <= 9'b1111010;
				8'b100001: c <= 9'b111000110;
				8'b1000110: c <= 9'b11111011;
				8'b1110010: c <= 9'b1010001;
				8'b1010000: c <= 9'b100110000;
				8'b1111010: c <= 9'b110001111;
				8'b1010101: c <= 9'b111001000;
				8'b111011: c <= 9'b101000110;
				8'b1001101: c <= 9'b11100111;
				8'b111111: c <= 9'b101010110;
				8'b1101110: c <= 9'b1;
				8'b1111011: c <= 9'b1000000;
				8'b1001011: c <= 9'b100101000;
				8'b1101111: c <= 9'b1010101;
				8'b1101000: c <= 9'b111101111;
				8'b101100: c <= 9'b111100111;
				8'b100100: c <= 9'b11101001;
				8'b1111000: c <= 9'b110111111;
				8'b1000101: c <= 9'b11001101;
				8'b1011001: c <= 9'b110010110;
				8'b110100: c <= 9'b111101111;
				8'b1111001: c <= 9'b110110011;
				8'b1110001: c <= 9'b10100100;
				8'b1001111: c <= 9'b1100;
				8'b1100101: c <= 9'b1101000;
				8'b1111110: c <= 9'b110101111;
				8'b1111100: c <= 9'b1100111;
				8'b1010110: c <= 9'b100110111;
				8'b110010: c <= 9'b1010111;
				8'b1101101: c <= 9'b101100101;
				8'b100011: c <= 9'b100011011;
				8'b1110101: c <= 9'b1110;
				8'b1111101: c <= 9'b101001101;
				8'b101001: c <= 9'b110011111;
				8'b1010010: c <= 9'b110001101;
				8'b1011000: c <= 9'b111101111;
				8'b101110: c <= 9'b101110111;
				8'b1000001: c <= 9'b1111011;
				default: c <= 9'b0;
			endcase
			9'b101001101 : case(di)
				8'b1000011: c <= 9'b110110101;
				8'b101000: c <= 9'b10011000;
				8'b111010: c <= 9'b111001100;
				8'b110110: c <= 9'b101100;
				8'b1100100: c <= 9'b101100011;
				8'b1000000: c <= 9'b1010110;
				8'b1110110: c <= 9'b100011111;
				8'b100101: c <= 9'b101100111;
				8'b101111: c <= 9'b1111010;
				8'b100110: c <= 9'b10100110;
				8'b1100011: c <= 9'b11011100;
				8'b1001000: c <= 9'b110111111;
				8'b111000: c <= 9'b100010000;
				8'b110001: c <= 9'b101100111;
				8'b1010111: c <= 9'b1100010;
				8'b1001110: c <= 9'b100101;
				8'b1101010: c <= 9'b110100110;
				8'b1001001: c <= 9'b100110110;
				8'b1100000: c <= 9'b10000001;
				8'b110111: c <= 9'b1010111;
				8'b1011101: c <= 9'b110100111;
				8'b1011011: c <= 9'b11110010;
				8'b111001: c <= 9'b1111111;
				8'b1001010: c <= 9'b100010100;
				8'b110011: c <= 9'b111111001;
				8'b1101100: c <= 9'b1100000;
				8'b1110111: c <= 9'b110100010;
				8'b101011: c <= 9'b111110101;
				8'b1101011: c <= 9'b101100011;
				8'b111100: c <= 9'b10011100;
				8'b1000111: c <= 9'b11000;
				8'b1011111: c <= 9'b10010;
				8'b1110100: c <= 9'b11111010;
				8'b101101: c <= 9'b100011010;
				8'b1010011: c <= 9'b101011;
				8'b1100001: c <= 9'b101110101;
				8'b110101: c <= 9'b101100010;
				8'b1000100: c <= 9'b1110111;
				8'b1010001: c <= 9'b10001011;
				8'b1010100: c <= 9'b111011010;
				8'b1100110: c <= 9'b101010101;
				8'b101010: c <= 9'b1000010;
				8'b1011110: c <= 9'b11011000;
				8'b1100111: c <= 9'b11100000;
				8'b1011010: c <= 9'b111101000;
				8'b1000010: c <= 9'b110011010;
				8'b111101: c <= 9'b11111000;
				8'b110000: c <= 9'b1101;
				8'b111110: c <= 9'b1001100;
				8'b1100010: c <= 9'b11011100;
				8'b1110000: c <= 9'b100011;
				8'b1101001: c <= 9'b110011000;
				8'b1110011: c <= 9'b100100110;
				8'b1001100: c <= 9'b11101000;
				8'b100001: c <= 9'b10101100;
				8'b1000110: c <= 9'b10000010;
				8'b1110010: c <= 9'b1001001;
				8'b1010000: c <= 9'b111000111;
				8'b1111010: c <= 9'b100000011;
				8'b1010101: c <= 9'b111001100;
				8'b111011: c <= 9'b101101000;
				8'b1001101: c <= 9'b101011000;
				8'b111111: c <= 9'b111110101;
				8'b1101110: c <= 9'b110100;
				8'b1111011: c <= 9'b11100100;
				8'b1001011: c <= 9'b101011111;
				8'b1101111: c <= 9'b111110101;
				8'b1101000: c <= 9'b100001010;
				8'b101100: c <= 9'b1100011;
				8'b100100: c <= 9'b101000110;
				8'b1111000: c <= 9'b111101;
				8'b1000101: c <= 9'b101100000;
				8'b1011001: c <= 9'b111011111;
				8'b110100: c <= 9'b1000001;
				8'b1111001: c <= 9'b101011;
				8'b1110001: c <= 9'b110100011;
				8'b1001111: c <= 9'b111101110;
				8'b1100101: c <= 9'b1111000;
				8'b1111110: c <= 9'b111010110;
				8'b1111100: c <= 9'b100000000;
				8'b1010110: c <= 9'b1101100;
				8'b110010: c <= 9'b11000010;
				8'b1101101: c <= 9'b11000000;
				8'b100011: c <= 9'b100000000;
				8'b1110101: c <= 9'b101101101;
				8'b1111101: c <= 9'b11111011;
				8'b101001: c <= 9'b111011100;
				8'b1010010: c <= 9'b100010110;
				8'b1011000: c <= 9'b11110111;
				8'b101110: c <= 9'b100010001;
				8'b1000001: c <= 9'b100111101;
				default: c <= 9'b0;
			endcase
			9'b11000001 : case(di)
				8'b1000011: c <= 9'b11;
				8'b101000: c <= 9'b101101001;
				8'b111010: c <= 9'b11111000;
				8'b110110: c <= 9'b10010011;
				8'b1100100: c <= 9'b101001011;
				8'b1000000: c <= 9'b11011101;
				8'b1110110: c <= 9'b111001101;
				8'b100101: c <= 9'b111010010;
				8'b101111: c <= 9'b111110110;
				8'b100110: c <= 9'b110100101;
				8'b1100011: c <= 9'b111000101;
				8'b1001000: c <= 9'b11110010;
				8'b111000: c <= 9'b11010011;
				8'b110001: c <= 9'b101010011;
				8'b1010111: c <= 9'b100011000;
				8'b1001110: c <= 9'b110000001;
				8'b1101010: c <= 9'b10001110;
				8'b1001001: c <= 9'b100010010;
				8'b1100000: c <= 9'b10100101;
				8'b110111: c <= 9'b110101101;
				8'b1011101: c <= 9'b101011000;
				8'b1011011: c <= 9'b10111000;
				8'b111001: c <= 9'b110010100;
				8'b1001010: c <= 9'b11010010;
				8'b110011: c <= 9'b10000011;
				8'b1101100: c <= 9'b101100101;
				8'b1110111: c <= 9'b111001000;
				8'b101011: c <= 9'b10100111;
				8'b1101011: c <= 9'b11111;
				8'b111100: c <= 9'b1111000;
				8'b1000111: c <= 9'b111100010;
				8'b1011111: c <= 9'b101010111;
				8'b1110100: c <= 9'b110110101;
				8'b101101: c <= 9'b101101;
				8'b1010011: c <= 9'b110110;
				8'b1100001: c <= 9'b110000001;
				8'b110101: c <= 9'b11110111;
				8'b1000100: c <= 9'b110110100;
				8'b1010001: c <= 9'b110000101;
				8'b1010100: c <= 9'b101110111;
				8'b1100110: c <= 9'b111111000;
				8'b101010: c <= 9'b10011;
				8'b1011110: c <= 9'b100010101;
				8'b1100111: c <= 9'b10011001;
				8'b1011010: c <= 9'b110111010;
				8'b1000010: c <= 9'b101111000;
				8'b111101: c <= 9'b10001110;
				8'b110000: c <= 9'b100000000;
				8'b111110: c <= 9'b1101110;
				8'b1100010: c <= 9'b10011011;
				8'b1110000: c <= 9'b110011100;
				8'b1101001: c <= 9'b101001;
				8'b1110011: c <= 9'b11011110;
				8'b1001100: c <= 9'b101101101;
				8'b100001: c <= 9'b101001100;
				8'b1000110: c <= 9'b100011001;
				8'b1110010: c <= 9'b111001011;
				8'b1010000: c <= 9'b11100011;
				8'b1111010: c <= 9'b10000011;
				8'b1010101: c <= 9'b100111010;
				8'b111011: c <= 9'b101100001;
				8'b1001101: c <= 9'b111111;
				8'b111111: c <= 9'b101101000;
				8'b1101110: c <= 9'b110001110;
				8'b1111011: c <= 9'b1101000;
				8'b1001011: c <= 9'b111001001;
				8'b1101111: c <= 9'b101110110;
				8'b1101000: c <= 9'b11111;
				8'b101100: c <= 9'b1000011;
				8'b100100: c <= 9'b100;
				8'b1111000: c <= 9'b11100010;
				8'b1000101: c <= 9'b110101011;
				8'b1011001: c <= 9'b10001110;
				8'b110100: c <= 9'b10011001;
				8'b1111001: c <= 9'b1000101;
				8'b1110001: c <= 9'b11111000;
				8'b1001111: c <= 9'b100001100;
				8'b1100101: c <= 9'b100011101;
				8'b1111110: c <= 9'b100001100;
				8'b1111100: c <= 9'b1001101;
				8'b1010110: c <= 9'b111100100;
				8'b110010: c <= 9'b110110;
				8'b1101101: c <= 9'b11010001;
				8'b100011: c <= 9'b111111001;
				8'b1110101: c <= 9'b1110111;
				8'b1111101: c <= 9'b10001111;
				8'b101001: c <= 9'b10101000;
				8'b1010010: c <= 9'b100001111;
				8'b1011000: c <= 9'b1101;
				8'b101110: c <= 9'b1111111;
				8'b1000001: c <= 9'b111110011;
				default: c <= 9'b0;
			endcase
			9'b11001 : case(di)
				8'b1000011: c <= 9'b110100001;
				8'b101000: c <= 9'b10010;
				8'b111010: c <= 9'b101100111;
				8'b110110: c <= 9'b111000;
				8'b1100100: c <= 9'b110111000;
				8'b1000000: c <= 9'b100011101;
				8'b1110110: c <= 9'b110011101;
				8'b100101: c <= 9'b10010110;
				8'b101111: c <= 9'b10111;
				8'b100110: c <= 9'b100110000;
				8'b1100011: c <= 9'b111100000;
				8'b1001000: c <= 9'b11100100;
				8'b111000: c <= 9'b1110000;
				8'b110001: c <= 9'b101100111;
				8'b1010111: c <= 9'b100111111;
				8'b1001110: c <= 9'b101110000;
				8'b1101010: c <= 9'b111101110;
				8'b1001001: c <= 9'b111101101;
				8'b1100000: c <= 9'b100101010;
				8'b110111: c <= 9'b101100100;
				8'b1011101: c <= 9'b101100101;
				8'b1011011: c <= 9'b10101;
				8'b111001: c <= 9'b111011101;
				8'b1001010: c <= 9'b100010110;
				8'b110011: c <= 9'b111001101;
				8'b1101100: c <= 9'b1011000;
				8'b1110111: c <= 9'b1000;
				8'b101011: c <= 9'b11001011;
				8'b1101011: c <= 9'b10000;
				8'b111100: c <= 9'b111011011;
				8'b1000111: c <= 9'b111001;
				8'b1011111: c <= 9'b101010;
				8'b1110100: c <= 9'b11100000;
				8'b101101: c <= 9'b110000101;
				8'b1010011: c <= 9'b10001100;
				8'b1100001: c <= 9'b100011010;
				8'b110101: c <= 9'b101101010;
				8'b1000100: c <= 9'b1010001;
				8'b1010001: c <= 9'b101110100;
				8'b1010100: c <= 9'b10010111;
				8'b1100110: c <= 9'b101000010;
				8'b101010: c <= 9'b1101101;
				8'b1011110: c <= 9'b110001010;
				8'b1100111: c <= 9'b1011100;
				8'b1011010: c <= 9'b111100111;
				8'b1000010: c <= 9'b1000111;
				8'b111101: c <= 9'b11001011;
				8'b110000: c <= 9'b111000;
				8'b111110: c <= 9'b10001110;
				8'b1100010: c <= 9'b10100110;
				8'b1110000: c <= 9'b1111100;
				8'b1101001: c <= 9'b10101100;
				8'b1110011: c <= 9'b1001101;
				8'b1001100: c <= 9'b111011001;
				8'b100001: c <= 9'b111010000;
				8'b1000110: c <= 9'b101001010;
				8'b1110010: c <= 9'b100000111;
				8'b1010000: c <= 9'b10101010;
				8'b1111010: c <= 9'b110110011;
				8'b1010101: c <= 9'b101011110;
				8'b111011: c <= 9'b10001110;
				8'b1001101: c <= 9'b11110010;
				8'b111111: c <= 9'b110100011;
				8'b1101110: c <= 9'b101101001;
				8'b1111011: c <= 9'b100101111;
				8'b1001011: c <= 9'b11110111;
				8'b1101111: c <= 9'b1001101;
				8'b1101000: c <= 9'b111010111;
				8'b101100: c <= 9'b110011;
				8'b100100: c <= 9'b11011100;
				8'b1111000: c <= 9'b100011000;
				8'b1000101: c <= 9'b111110001;
				8'b1011001: c <= 9'b100101110;
				8'b110100: c <= 9'b11100110;
				8'b1111001: c <= 9'b100100001;
				8'b1110001: c <= 9'b10111111;
				8'b1001111: c <= 9'b110011111;
				8'b1100101: c <= 9'b1101;
				8'b1111110: c <= 9'b11011000;
				8'b1111100: c <= 9'b111011010;
				8'b1010110: c <= 9'b111001111;
				8'b110010: c <= 9'b1101111;
				8'b1101101: c <= 9'b110100011;
				8'b100011: c <= 9'b101011011;
				8'b1110101: c <= 9'b110001001;
				8'b1111101: c <= 9'b111101000;
				8'b101001: c <= 9'b100100011;
				8'b1010010: c <= 9'b10011100;
				8'b1011000: c <= 9'b110000;
				8'b101110: c <= 9'b101001011;
				8'b1000001: c <= 9'b101000011;
				default: c <= 9'b0;
			endcase
			9'b100101111 : case(di)
				8'b1000011: c <= 9'b1111101;
				8'b101000: c <= 9'b100110110;
				8'b111010: c <= 9'b10000101;
				8'b110110: c <= 9'b11110110;
				8'b1100100: c <= 9'b100000001;
				8'b1000000: c <= 9'b110110010;
				8'b1110110: c <= 9'b1110;
				8'b100101: c <= 9'b101011011;
				8'b101111: c <= 9'b100100010;
				8'b100110: c <= 9'b100011011;
				8'b1100011: c <= 9'b10011001;
				8'b1001000: c <= 9'b10011010;
				8'b111000: c <= 9'b11001010;
				8'b110001: c <= 9'b111000000;
				8'b1010111: c <= 9'b11111110;
				8'b1001110: c <= 9'b1001;
				8'b1101010: c <= 9'b110011110;
				8'b1001001: c <= 9'b101000100;
				8'b1100000: c <= 9'b11011000;
				8'b110111: c <= 9'b11101111;
				8'b1011101: c <= 9'b111001110;
				8'b1011011: c <= 9'b11011011;
				8'b111001: c <= 9'b1000101;
				8'b1001010: c <= 9'b100001;
				8'b110011: c <= 9'b111;
				8'b1101100: c <= 9'b100001110;
				8'b1110111: c <= 9'b110010011;
				8'b101011: c <= 9'b110011001;
				8'b1101011: c <= 9'b11101101;
				8'b111100: c <= 9'b11101011;
				8'b1000111: c <= 9'b10101000;
				8'b1011111: c <= 9'b100010010;
				8'b1110100: c <= 9'b10011011;
				8'b101101: c <= 9'b110110101;
				8'b1010011: c <= 9'b110001001;
				8'b1100001: c <= 9'b10111100;
				8'b110101: c <= 9'b111000010;
				8'b1000100: c <= 9'b1000010;
				8'b1010001: c <= 9'b10100;
				8'b1010100: c <= 9'b110000111;
				8'b1100110: c <= 9'b1;
				8'b101010: c <= 9'b100001001;
				8'b1011110: c <= 9'b1110011;
				8'b1100111: c <= 9'b100110000;
				8'b1011010: c <= 9'b111101111;
				8'b1000010: c <= 9'b1100011;
				8'b111101: c <= 9'b100000000;
				8'b110000: c <= 9'b11000;
				8'b111110: c <= 9'b101111000;
				8'b1100010: c <= 9'b10100101;
				8'b1110000: c <= 9'b1011110;
				8'b1101001: c <= 9'b111110001;
				8'b1110011: c <= 9'b111101;
				8'b1001100: c <= 9'b101110000;
				8'b100001: c <= 9'b110001100;
				8'b1000110: c <= 9'b111100000;
				8'b1110010: c <= 9'b1001101;
				8'b1010000: c <= 9'b1110001;
				8'b1111010: c <= 9'b111101100;
				8'b1010101: c <= 9'b10111101;
				8'b111011: c <= 9'b111010111;
				8'b1001101: c <= 9'b111001010;
				8'b111111: c <= 9'b100110010;
				8'b1101110: c <= 9'b111001;
				8'b1111011: c <= 9'b100010011;
				8'b1001011: c <= 9'b100010011;
				8'b1101111: c <= 9'b10010101;
				8'b1101000: c <= 9'b10011100;
				8'b101100: c <= 9'b101011110;
				8'b100100: c <= 9'b101010010;
				8'b1111000: c <= 9'b101110110;
				8'b1000101: c <= 9'b100000100;
				8'b1011001: c <= 9'b1101110;
				8'b110100: c <= 9'b111;
				8'b1111001: c <= 9'b111100110;
				8'b1110001: c <= 9'b1011010;
				8'b1001111: c <= 9'b11001000;
				8'b1100101: c <= 9'b10011000;
				8'b1111110: c <= 9'b111001010;
				8'b1111100: c <= 9'b110011111;
				8'b1010110: c <= 9'b100100111;
				8'b110010: c <= 9'b111011111;
				8'b1101101: c <= 9'b100001111;
				8'b100011: c <= 9'b11001110;
				8'b1110101: c <= 9'b1000111;
				8'b1111101: c <= 9'b10001000;
				8'b101001: c <= 9'b11011001;
				8'b1010010: c <= 9'b1100110;
				8'b1011000: c <= 9'b10001111;
				8'b101110: c <= 9'b111001;
				8'b1000001: c <= 9'b100011011;
				default: c <= 9'b0;
			endcase
			9'b11 : case(di)
				8'b1000011: c <= 9'b11100000;
				8'b101000: c <= 9'b111101001;
				8'b111010: c <= 9'b101101010;
				8'b110110: c <= 9'b1110101;
				8'b1100100: c <= 9'b100100000;
				8'b1000000: c <= 9'b10110110;
				8'b1110110: c <= 9'b10010101;
				8'b100101: c <= 9'b100111111;
				8'b101111: c <= 9'b101000010;
				8'b100110: c <= 9'b10000;
				8'b1100011: c <= 9'b111101000;
				8'b1001000: c <= 9'b11100000;
				8'b111000: c <= 9'b110;
				8'b110001: c <= 9'b110010010;
				8'b1010111: c <= 9'b111011100;
				8'b1001110: c <= 9'b100100;
				8'b1101010: c <= 9'b111111011;
				8'b1001001: c <= 9'b10010;
				8'b1100000: c <= 9'b110110100;
				8'b110111: c <= 9'b11000;
				8'b1011101: c <= 9'b11100100;
				8'b1011011: c <= 9'b11101100;
				8'b111001: c <= 9'b100100001;
				8'b1001010: c <= 9'b110001001;
				8'b110011: c <= 9'b110011100;
				8'b1101100: c <= 9'b10101011;
				8'b1110111: c <= 9'b11110010;
				8'b101011: c <= 9'b111101001;
				8'b1101011: c <= 9'b100000100;
				8'b111100: c <= 9'b100000011;
				8'b1000111: c <= 9'b11101011;
				8'b1011111: c <= 9'b100110101;
				8'b1110100: c <= 9'b111110000;
				8'b101101: c <= 9'b1011000;
				8'b1010011: c <= 9'b110011110;
				8'b1100001: c <= 9'b101101010;
				8'b110101: c <= 9'b110111011;
				8'b1000100: c <= 9'b111111;
				8'b1010001: c <= 9'b11110010;
				8'b1010100: c <= 9'b111000100;
				8'b1100110: c <= 9'b101011011;
				8'b101010: c <= 9'b10111010;
				8'b1011110: c <= 9'b1010000;
				8'b1100111: c <= 9'b11101;
				8'b1011010: c <= 9'b1101110;
				8'b1000010: c <= 9'b111011100;
				8'b111101: c <= 9'b100111100;
				8'b110000: c <= 9'b110101011;
				8'b111110: c <= 9'b1110000;
				8'b1100010: c <= 9'b101100011;
				8'b1110000: c <= 9'b101001011;
				8'b1101001: c <= 9'b110110011;
				8'b1110011: c <= 9'b11110000;
				8'b1001100: c <= 9'b100011000;
				8'b100001: c <= 9'b11101111;
				8'b1000110: c <= 9'b1100101;
				8'b1110010: c <= 9'b1010001;
				8'b1010000: c <= 9'b10110100;
				8'b1111010: c <= 9'b100001011;
				8'b1010101: c <= 9'b110010010;
				8'b111011: c <= 9'b111010000;
				8'b1001101: c <= 9'b11110110;
				8'b111111: c <= 9'b101100;
				8'b1101110: c <= 9'b111;
				8'b1111011: c <= 9'b100101010;
				8'b1001011: c <= 9'b101000101;
				8'b1101111: c <= 9'b101010011;
				8'b1101000: c <= 9'b110010110;
				8'b101100: c <= 9'b1111011;
				8'b100100: c <= 9'b111111110;
				8'b1111000: c <= 9'b1011100;
				8'b1000101: c <= 9'b11010000;
				8'b1011001: c <= 9'b110111100;
				8'b110100: c <= 9'b110101111;
				8'b1111001: c <= 9'b110110000;
				8'b1110001: c <= 9'b10010;
				8'b1001111: c <= 9'b100010010;
				8'b1100101: c <= 9'b101010000;
				8'b1111110: c <= 9'b11001101;
				8'b1111100: c <= 9'b10000010;
				8'b1010110: c <= 9'b110110011;
				8'b110010: c <= 9'b110111001;
				8'b1101101: c <= 9'b110100010;
				8'b100011: c <= 9'b1000111;
				8'b1110101: c <= 9'b101110111;
				8'b1111101: c <= 9'b1111000;
				8'b101001: c <= 9'b1111000;
				8'b1010010: c <= 9'b101110010;
				8'b1011000: c <= 9'b10101101;
				8'b101110: c <= 9'b10110100;
				8'b1000001: c <= 9'b101001110;
				default: c <= 9'b0;
			endcase
			9'b100010110 : case(di)
				8'b1000011: c <= 9'b100011101;
				8'b101000: c <= 9'b1000100;
				8'b111010: c <= 9'b101010000;
				8'b110110: c <= 9'b110110010;
				8'b1100100: c <= 9'b11000100;
				8'b1000000: c <= 9'b110000010;
				8'b1110110: c <= 9'b1001011;
				8'b100101: c <= 9'b111011;
				8'b101111: c <= 9'b101111000;
				8'b100110: c <= 9'b1011001;
				8'b1100011: c <= 9'b111111101;
				8'b1001000: c <= 9'b11001110;
				8'b111000: c <= 9'b11010011;
				8'b110001: c <= 9'b111000101;
				8'b1010111: c <= 9'b100001011;
				8'b1001110: c <= 9'b10001110;
				8'b1101010: c <= 9'b110111001;
				8'b1001001: c <= 9'b100001001;
				8'b1100000: c <= 9'b100100001;
				8'b110111: c <= 9'b101101000;
				8'b1011101: c <= 9'b10100110;
				8'b1011011: c <= 9'b11110000;
				8'b111001: c <= 9'b100101000;
				8'b1001010: c <= 9'b10111000;
				8'b110011: c <= 9'b110011110;
				8'b1101100: c <= 9'b110010100;
				8'b1110111: c <= 9'b10101110;
				8'b101011: c <= 9'b100010011;
				8'b1101011: c <= 9'b11;
				8'b111100: c <= 9'b101100110;
				8'b1000111: c <= 9'b10111010;
				8'b1011111: c <= 9'b110010101;
				8'b1110100: c <= 9'b100101010;
				8'b101101: c <= 9'b110010;
				8'b1010011: c <= 9'b11001010;
				8'b1100001: c <= 9'b111111;
				8'b110101: c <= 9'b11000100;
				8'b1000100: c <= 9'b101101001;
				8'b1010001: c <= 9'b11011;
				8'b1010100: c <= 9'b100100010;
				8'b1100110: c <= 9'b11001001;
				8'b101010: c <= 9'b111001;
				8'b1011110: c <= 9'b111010100;
				8'b1100111: c <= 9'b10011100;
				8'b1011010: c <= 9'b111110000;
				8'b1000010: c <= 9'b10111110;
				8'b111101: c <= 9'b1101;
				8'b110000: c <= 9'b110011001;
				8'b111110: c <= 9'b1111110;
				8'b1100010: c <= 9'b1011000;
				8'b1110000: c <= 9'b100000101;
				8'b1101001: c <= 9'b10101101;
				8'b1110011: c <= 9'b11100100;
				8'b1001100: c <= 9'b10110111;
				8'b100001: c <= 9'b11010011;
				8'b1000110: c <= 9'b100111111;
				8'b1110010: c <= 9'b10011101;
				8'b1010000: c <= 9'b110001010;
				8'b1111010: c <= 9'b110001;
				8'b1010101: c <= 9'b100111110;
				8'b111011: c <= 9'b101101111;
				8'b1001101: c <= 9'b10100111;
				8'b111111: c <= 9'b10100101;
				8'b1101110: c <= 9'b111111011;
				8'b1111011: c <= 9'b101011110;
				8'b1001011: c <= 9'b1001101;
				8'b1101111: c <= 9'b111010100;
				8'b1101000: c <= 9'b1000;
				8'b101100: c <= 9'b110101;
				8'b100100: c <= 9'b100001100;
				8'b1111000: c <= 9'b11000110;
				8'b1000101: c <= 9'b101000011;
				8'b1011001: c <= 9'b1101000;
				8'b110100: c <= 9'b101000;
				8'b1111001: c <= 9'b101000001;
				8'b1110001: c <= 9'b1100000;
				8'b1001111: c <= 9'b100010100;
				8'b1100101: c <= 9'b100001001;
				8'b1111110: c <= 9'b10000110;
				8'b1111100: c <= 9'b110000011;
				8'b1010110: c <= 9'b11001110;
				8'b110010: c <= 9'b100101100;
				8'b1101101: c <= 9'b110001101;
				8'b100011: c <= 9'b100001011;
				8'b1110101: c <= 9'b10100101;
				8'b1111101: c <= 9'b111011;
				8'b101001: c <= 9'b1000101;
				8'b1010010: c <= 9'b1001101;
				8'b1011000: c <= 9'b101110011;
				8'b101110: c <= 9'b100111101;
				8'b1000001: c <= 9'b11111010;
				default: c <= 9'b0;
			endcase
			9'b10101111 : case(di)
				8'b1000011: c <= 9'b101101100;
				8'b101000: c <= 9'b101110010;
				8'b111010: c <= 9'b110111110;
				8'b110110: c <= 9'b110101010;
				8'b1100100: c <= 9'b101010110;
				8'b1000000: c <= 9'b1001000;
				8'b1110110: c <= 9'b1100111;
				8'b100101: c <= 9'b100101011;
				8'b101111: c <= 9'b11111000;
				8'b100110: c <= 9'b101011010;
				8'b1100011: c <= 9'b100000000;
				8'b1001000: c <= 9'b110100000;
				8'b111000: c <= 9'b110011100;
				8'b110001: c <= 9'b1001001;
				8'b1010111: c <= 9'b101101011;
				8'b1001110: c <= 9'b110100;
				8'b1101010: c <= 9'b101101011;
				8'b1001001: c <= 9'b101101;
				8'b1100000: c <= 9'b10001000;
				8'b110111: c <= 9'b1100;
				8'b1011101: c <= 9'b101010101;
				8'b1011011: c <= 9'b101110101;
				8'b111001: c <= 9'b110111111;
				8'b1001010: c <= 9'b100001;
				8'b110011: c <= 9'b100001001;
				8'b1101100: c <= 9'b100100111;
				8'b1110111: c <= 9'b101101000;
				8'b101011: c <= 9'b110100010;
				8'b1101011: c <= 9'b111111;
				8'b111100: c <= 9'b100111001;
				8'b1000111: c <= 9'b111001001;
				8'b1011111: c <= 9'b1111111;
				8'b1110100: c <= 9'b110111110;
				8'b101101: c <= 9'b101110;
				8'b1010011: c <= 9'b101010;
				8'b1100001: c <= 9'b101110100;
				8'b110101: c <= 9'b110001011;
				8'b1000100: c <= 9'b110111110;
				8'b1010001: c <= 9'b110010111;
				8'b1010100: c <= 9'b100000011;
				8'b1100110: c <= 9'b10010;
				8'b101010: c <= 9'b100110010;
				8'b1011110: c <= 9'b1011010;
				8'b1100111: c <= 9'b111101110;
				8'b1011010: c <= 9'b111111110;
				8'b1000010: c <= 9'b101110000;
				8'b111101: c <= 9'b1101010;
				8'b110000: c <= 9'b111111111;
				8'b111110: c <= 9'b10100100;
				8'b1100010: c <= 9'b101010111;
				8'b1110000: c <= 9'b1111111;
				8'b1101001: c <= 9'b111001010;
				8'b1110011: c <= 9'b110;
				8'b1001100: c <= 9'b111110101;
				8'b100001: c <= 9'b100000110;
				8'b1000110: c <= 9'b11110101;
				8'b1110010: c <= 9'b10011111;
				8'b1010000: c <= 9'b101100010;
				8'b1111010: c <= 9'b110011011;
				8'b1010101: c <= 9'b1000;
				8'b111011: c <= 9'b110101110;
				8'b1001101: c <= 9'b11010111;
				8'b111111: c <= 9'b111100;
				8'b1101110: c <= 9'b11000110;
				8'b1111011: c <= 9'b101010001;
				8'b1001011: c <= 9'b101010111;
				8'b1101111: c <= 9'b111011101;
				8'b1101000: c <= 9'b11000100;
				8'b101100: c <= 9'b100011011;
				8'b100100: c <= 9'b111000101;
				8'b1111000: c <= 9'b11111011;
				8'b1000101: c <= 9'b111000011;
				8'b1011001: c <= 9'b111101111;
				8'b110100: c <= 9'b101000111;
				8'b1111001: c <= 9'b1001111;
				8'b1110001: c <= 9'b111011011;
				8'b1001111: c <= 9'b10111000;
				8'b1100101: c <= 9'b101100100;
				8'b1111110: c <= 9'b110100010;
				8'b1111100: c <= 9'b11001111;
				8'b1010110: c <= 9'b100001111;
				8'b110010: c <= 9'b101000001;
				8'b1101101: c <= 9'b10111111;
				8'b100011: c <= 9'b1100101;
				8'b1110101: c <= 9'b10110100;
				8'b1111101: c <= 9'b100010010;
				8'b101001: c <= 9'b111111;
				8'b1010010: c <= 9'b1011011;
				8'b1011000: c <= 9'b111111;
				8'b101110: c <= 9'b101011010;
				8'b1000001: c <= 9'b1001101;
				default: c <= 9'b0;
			endcase
			9'b111001001 : case(di)
				8'b1000011: c <= 9'b100100000;
				8'b101000: c <= 9'b111100111;
				8'b111010: c <= 9'b111011001;
				8'b110110: c <= 9'b101011101;
				8'b1100100: c <= 9'b111011110;
				8'b1000000: c <= 9'b1100101;
				8'b1110110: c <= 9'b101100100;
				8'b100101: c <= 9'b10100011;
				8'b101111: c <= 9'b110101001;
				8'b100110: c <= 9'b101011;
				8'b1100011: c <= 9'b10111000;
				8'b1001000: c <= 9'b10000010;
				8'b111000: c <= 9'b111101;
				8'b110001: c <= 9'b10001010;
				8'b1010111: c <= 9'b11100111;
				8'b1001110: c <= 9'b100000110;
				8'b1101010: c <= 9'b111000110;
				8'b1001001: c <= 9'b10010110;
				8'b1100000: c <= 9'b1110011;
				8'b110111: c <= 9'b111111111;
				8'b1011101: c <= 9'b111011;
				8'b1011011: c <= 9'b10011;
				8'b111001: c <= 9'b10101110;
				8'b1001010: c <= 9'b100101;
				8'b110011: c <= 9'b101001100;
				8'b1101100: c <= 9'b111001100;
				8'b1110111: c <= 9'b10011011;
				8'b101011: c <= 9'b101000110;
				8'b1101011: c <= 9'b1000110;
				8'b111100: c <= 9'b110001011;
				8'b1000111: c <= 9'b1110111;
				8'b1011111: c <= 9'b100101101;
				8'b1110100: c <= 9'b110110110;
				8'b101101: c <= 9'b10111101;
				8'b1010011: c <= 9'b111000100;
				8'b1100001: c <= 9'b10010111;
				8'b110101: c <= 9'b101001111;
				8'b1000100: c <= 9'b11001101;
				8'b1010001: c <= 9'b101011101;
				8'b1010100: c <= 9'b110000110;
				8'b1100110: c <= 9'b101011001;
				8'b101010: c <= 9'b11001111;
				8'b1011110: c <= 9'b11010100;
				8'b1100111: c <= 9'b11100100;
				8'b1011010: c <= 9'b11001001;
				8'b1000010: c <= 9'b111100100;
				8'b111101: c <= 9'b1101001;
				8'b110000: c <= 9'b111101110;
				8'b111110: c <= 9'b111101110;
				8'b1100010: c <= 9'b111100001;
				8'b1110000: c <= 9'b11010011;
				8'b1101001: c <= 9'b10010000;
				8'b1110011: c <= 9'b111000100;
				8'b1001100: c <= 9'b100010111;
				8'b100001: c <= 9'b1100100;
				8'b1000110: c <= 9'b100100110;
				8'b1110010: c <= 9'b110101;
				8'b1010000: c <= 9'b101100111;
				8'b1111010: c <= 9'b1111110;
				8'b1010101: c <= 9'b10000000;
				8'b111011: c <= 9'b111101000;
				8'b1001101: c <= 9'b1110000;
				8'b111111: c <= 9'b111111;
				8'b1101110: c <= 9'b11100111;
				8'b1111011: c <= 9'b110011011;
				8'b1001011: c <= 9'b111110000;
				8'b1101111: c <= 9'b101110011;
				8'b1101000: c <= 9'b10101000;
				8'b101100: c <= 9'b111101000;
				8'b100100: c <= 9'b111101110;
				8'b1111000: c <= 9'b11001110;
				8'b1000101: c <= 9'b10001000;
				8'b1011001: c <= 9'b111101100;
				8'b110100: c <= 9'b11111101;
				8'b1111001: c <= 9'b10100100;
				8'b1110001: c <= 9'b10101011;
				8'b1001111: c <= 9'b101010;
				8'b1100101: c <= 9'b111100110;
				8'b1111110: c <= 9'b11011000;
				8'b1111100: c <= 9'b1000110;
				8'b1010110: c <= 9'b100011001;
				8'b110010: c <= 9'b100110101;
				8'b1101101: c <= 9'b1100101;
				8'b100011: c <= 9'b1101;
				8'b1110101: c <= 9'b110010;
				8'b1111101: c <= 9'b11110001;
				8'b101001: c <= 9'b11111;
				8'b1010010: c <= 9'b110100110;
				8'b1011000: c <= 9'b111001000;
				8'b101110: c <= 9'b10101011;
				8'b1000001: c <= 9'b10101011;
				default: c <= 9'b0;
			endcase
			9'b110100 : case(di)
				8'b1000011: c <= 9'b1111;
				8'b101000: c <= 9'b1010001;
				8'b111010: c <= 9'b100100000;
				8'b110110: c <= 9'b1111100;
				8'b1100100: c <= 9'b111000100;
				8'b1000000: c <= 9'b10111101;
				8'b1110110: c <= 9'b10101010;
				8'b100101: c <= 9'b1000110;
				8'b101111: c <= 9'b1110011;
				8'b100110: c <= 9'b10000111;
				8'b1100011: c <= 9'b1000100;
				8'b1001000: c <= 9'b100101101;
				8'b111000: c <= 9'b101001001;
				8'b110001: c <= 9'b110111100;
				8'b1010111: c <= 9'b101100001;
				8'b1001110: c <= 9'b101100111;
				8'b1101010: c <= 9'b11010111;
				8'b1001001: c <= 9'b110010111;
				8'b1100000: c <= 9'b111110000;
				8'b110111: c <= 9'b11011001;
				8'b1011101: c <= 9'b110110000;
				8'b1011011: c <= 9'b100111100;
				8'b111001: c <= 9'b11100010;
				8'b1001010: c <= 9'b101010101;
				8'b110011: c <= 9'b101110011;
				8'b1101100: c <= 9'b1110100;
				8'b1110111: c <= 9'b110100010;
				8'b101011: c <= 9'b1101111;
				8'b1101011: c <= 9'b111010100;
				8'b111100: c <= 9'b10110101;
				8'b1000111: c <= 9'b100101101;
				8'b1011111: c <= 9'b101110011;
				8'b1110100: c <= 9'b110101111;
				8'b101101: c <= 9'b110000111;
				8'b1010011: c <= 9'b1011001;
				8'b1100001: c <= 9'b10100000;
				8'b110101: c <= 9'b100010111;
				8'b1000100: c <= 9'b111100011;
				8'b1010001: c <= 9'b11100010;
				8'b1010100: c <= 9'b1110010;
				8'b1100110: c <= 9'b11110010;
				8'b101010: c <= 9'b111010100;
				8'b1011110: c <= 9'b100010111;
				8'b1100111: c <= 9'b100000011;
				8'b1011010: c <= 9'b111100100;
				8'b1000010: c <= 9'b101000011;
				8'b111101: c <= 9'b11111000;
				8'b110000: c <= 9'b11000;
				8'b111110: c <= 9'b110011110;
				8'b1100010: c <= 9'b100001101;
				8'b1110000: c <= 9'b1111101;
				8'b1101001: c <= 9'b10100;
				8'b1110011: c <= 9'b1111010;
				8'b1001100: c <= 9'b111001011;
				8'b100001: c <= 9'b100001;
				8'b1000110: c <= 9'b111101001;
				8'b1110010: c <= 9'b110111111;
				8'b1010000: c <= 9'b100001111;
				8'b1111010: c <= 9'b111110001;
				8'b1010101: c <= 9'b110101100;
				8'b111011: c <= 9'b101000011;
				8'b1001101: c <= 9'b101000001;
				8'b111111: c <= 9'b110111;
				8'b1101110: c <= 9'b10011011;
				8'b1111011: c <= 9'b11011100;
				8'b1001011: c <= 9'b111111000;
				8'b1101111: c <= 9'b110000111;
				8'b1101000: c <= 9'b11100110;
				8'b101100: c <= 9'b111001010;
				8'b100100: c <= 9'b111101111;
				8'b1111000: c <= 9'b101101110;
				8'b1000101: c <= 9'b10111100;
				8'b1011001: c <= 9'b101101001;
				8'b110100: c <= 9'b1110000;
				8'b1111001: c <= 9'b101010110;
				8'b1110001: c <= 9'b10110111;
				8'b1001111: c <= 9'b110001011;
				8'b1100101: c <= 9'b10100101;
				8'b1111110: c <= 9'b111100000;
				8'b1111100: c <= 9'b10011;
				8'b1010110: c <= 9'b101001000;
				8'b110010: c <= 9'b110011101;
				8'b1101101: c <= 9'b100111001;
				8'b100011: c <= 9'b110100;
				8'b1110101: c <= 9'b10111010;
				8'b1111101: c <= 9'b100001100;
				8'b101001: c <= 9'b111001101;
				8'b1010010: c <= 9'b10111001;
				8'b1011000: c <= 9'b101111010;
				8'b101110: c <= 9'b110011101;
				8'b1000001: c <= 9'b101010000;
				default: c <= 9'b0;
			endcase
			9'b1000 : case(di)
				8'b1000011: c <= 9'b10000111;
				8'b101000: c <= 9'b101101101;
				8'b111010: c <= 9'b100111000;
				8'b110110: c <= 9'b11011001;
				8'b1100100: c <= 9'b101010101;
				8'b1000000: c <= 9'b101110110;
				8'b1110110: c <= 9'b110100011;
				8'b100101: c <= 9'b110000;
				8'b101111: c <= 9'b110100000;
				8'b100110: c <= 9'b1110010;
				8'b1100011: c <= 9'b110100;
				8'b1001000: c <= 9'b110110010;
				8'b111000: c <= 9'b10111110;
				8'b110001: c <= 9'b110011001;
				8'b1010111: c <= 9'b11011;
				8'b1001110: c <= 9'b1111001;
				8'b1101010: c <= 9'b101101001;
				8'b1001001: c <= 9'b111111;
				8'b1100000: c <= 9'b101000100;
				8'b110111: c <= 9'b111010110;
				8'b1011101: c <= 9'b101111010;
				8'b1011011: c <= 9'b111110110;
				8'b111001: c <= 9'b100110101;
				8'b1001010: c <= 9'b100001100;
				8'b110011: c <= 9'b10101100;
				8'b1101100: c <= 9'b10000111;
				8'b1110111: c <= 9'b1110001;
				8'b101011: c <= 9'b11101100;
				8'b1101011: c <= 9'b100000000;
				8'b111100: c <= 9'b100010111;
				8'b1000111: c <= 9'b1100101;
				8'b1011111: c <= 9'b11110000;
				8'b1110100: c <= 9'b11000010;
				8'b101101: c <= 9'b110010101;
				8'b1010011: c <= 9'b111010110;
				8'b1100001: c <= 9'b100110110;
				8'b110101: c <= 9'b100010110;
				8'b1000100: c <= 9'b1111011;
				8'b1010001: c <= 9'b111111000;
				8'b1010100: c <= 9'b111110011;
				8'b1100110: c <= 9'b11000001;
				8'b101010: c <= 9'b110101001;
				8'b1011110: c <= 9'b111101101;
				8'b1100111: c <= 9'b101101001;
				8'b1011010: c <= 9'b110000010;
				8'b1000010: c <= 9'b100110110;
				8'b111101: c <= 9'b11111001;
				8'b110000: c <= 9'b1010000;
				8'b111110: c <= 9'b11100110;
				8'b1100010: c <= 9'b100011;
				8'b1110000: c <= 9'b11001101;
				8'b1101001: c <= 9'b100101011;
				8'b1110011: c <= 9'b100100000;
				8'b1001100: c <= 9'b11111101;
				8'b100001: c <= 9'b101110111;
				8'b1000110: c <= 9'b101001100;
				8'b1110010: c <= 9'b1110100;
				8'b1010000: c <= 9'b110111010;
				8'b1111010: c <= 9'b100101000;
				8'b1010101: c <= 9'b100101111;
				8'b111011: c <= 9'b10001010;
				8'b1001101: c <= 9'b110011001;
				8'b111111: c <= 9'b101100001;
				8'b1101110: c <= 9'b101010011;
				8'b1111011: c <= 9'b100101001;
				8'b1001011: c <= 9'b101110011;
				8'b1101111: c <= 9'b110100110;
				8'b1101000: c <= 9'b11111110;
				8'b101100: c <= 9'b1101101;
				8'b100100: c <= 9'b10111011;
				8'b1111000: c <= 9'b11011000;
				8'b1000101: c <= 9'b11001011;
				8'b1011001: c <= 9'b1100111;
				8'b110100: c <= 9'b110011000;
				8'b1111001: c <= 9'b110001010;
				8'b1110001: c <= 9'b11110101;
				8'b1001111: c <= 9'b101000;
				8'b1100101: c <= 9'b111011;
				8'b1111110: c <= 9'b101100001;
				8'b1111100: c <= 9'b110111100;
				8'b1010110: c <= 9'b111110001;
				8'b110010: c <= 9'b10110110;
				8'b1101101: c <= 9'b101011111;
				8'b100011: c <= 9'b100111110;
				8'b1110101: c <= 9'b111100100;
				8'b1111101: c <= 9'b1101110;
				8'b101001: c <= 9'b10110101;
				8'b1010010: c <= 9'b1010011;
				8'b1011000: c <= 9'b100000110;
				8'b101110: c <= 9'b11111010;
				8'b1000001: c <= 9'b111000000;
				default: c <= 9'b0;
			endcase
			9'b11100001 : case(di)
				8'b1000011: c <= 9'b10001011;
				8'b101000: c <= 9'b100101011;
				8'b111010: c <= 9'b1001;
				8'b110110: c <= 9'b110111001;
				8'b1100100: c <= 9'b110000011;
				8'b1000000: c <= 9'b111011;
				8'b1110110: c <= 9'b101011001;
				8'b100101: c <= 9'b110111010;
				8'b101111: c <= 9'b11100001;
				8'b100110: c <= 9'b101101011;
				8'b1100011: c <= 9'b100010000;
				8'b1001000: c <= 9'b111101000;
				8'b111000: c <= 9'b10001101;
				8'b110001: c <= 9'b101001001;
				8'b1010111: c <= 9'b101110100;
				8'b1001110: c <= 9'b101010100;
				8'b1101010: c <= 9'b110110111;
				8'b1001001: c <= 9'b111000011;
				8'b1100000: c <= 9'b100001110;
				8'b110111: c <= 9'b10001100;
				8'b1011101: c <= 9'b11010011;
				8'b1011011: c <= 9'b1101010;
				8'b111001: c <= 9'b100101010;
				8'b1001010: c <= 9'b111110101;
				8'b110011: c <= 9'b101111001;
				8'b1101100: c <= 9'b10110100;
				8'b1110111: c <= 9'b10111000;
				8'b101011: c <= 9'b11100011;
				8'b1101011: c <= 9'b101100110;
				8'b111100: c <= 9'b111111010;
				8'b1000111: c <= 9'b10100110;
				8'b1011111: c <= 9'b11;
				8'b1110100: c <= 9'b1110001;
				8'b101101: c <= 9'b100110110;
				8'b1010011: c <= 9'b11001001;
				8'b1100001: c <= 9'b101001010;
				8'b110101: c <= 9'b1101100;
				8'b1000100: c <= 9'b111011010;
				8'b1010001: c <= 9'b110011110;
				8'b1010100: c <= 9'b111111001;
				8'b1100110: c <= 9'b1010011;
				8'b101010: c <= 9'b1110111;
				8'b1011110: c <= 9'b100101110;
				8'b1100111: c <= 9'b100010110;
				8'b1011010: c <= 9'b110000000;
				8'b1000010: c <= 9'b10000001;
				8'b111101: c <= 9'b101000010;
				8'b110000: c <= 9'b1011111;
				8'b111110: c <= 9'b1110101;
				8'b1100010: c <= 9'b10001101;
				8'b1110000: c <= 9'b10010;
				8'b1101001: c <= 9'b110010110;
				8'b1110011: c <= 9'b100010001;
				8'b1001100: c <= 9'b11100;
				8'b100001: c <= 9'b100000000;
				8'b1000110: c <= 9'b101100000;
				8'b1110010: c <= 9'b1010111;
				8'b1010000: c <= 9'b10111011;
				8'b1111010: c <= 9'b101001100;
				8'b1010101: c <= 9'b1010111;
				8'b111011: c <= 9'b111111111;
				8'b1001101: c <= 9'b101110111;
				8'b111111: c <= 9'b11100001;
				8'b1101110: c <= 9'b110100000;
				8'b1111011: c <= 9'b100101011;
				8'b1001011: c <= 9'b111001100;
				8'b1101111: c <= 9'b1110001;
				8'b1101000: c <= 9'b101100100;
				8'b101100: c <= 9'b11110111;
				8'b100100: c <= 9'b101110001;
				8'b1111000: c <= 9'b101110001;
				8'b1000101: c <= 9'b110001110;
				8'b1011001: c <= 9'b101000111;
				8'b110100: c <= 9'b1101;
				8'b1111001: c <= 9'b110111010;
				8'b1110001: c <= 9'b1110111;
				8'b1001111: c <= 9'b101100101;
				8'b1100101: c <= 9'b101100101;
				8'b1111110: c <= 9'b10001100;
				8'b1111100: c <= 9'b1111101;
				8'b1010110: c <= 9'b1011010;
				8'b110010: c <= 9'b11010;
				8'b1101101: c <= 9'b1011110;
				8'b100011: c <= 9'b100100011;
				8'b1110101: c <= 9'b10111000;
				8'b1111101: c <= 9'b10100;
				8'b101001: c <= 9'b111000000;
				8'b1010010: c <= 9'b100101001;
				8'b1011000: c <= 9'b110010;
				8'b101110: c <= 9'b101100010;
				8'b1000001: c <= 9'b11011101;
				default: c <= 9'b0;
			endcase
			9'b111111110 : case(di)
				8'b1000011: c <= 9'b111011110;
				8'b101000: c <= 9'b100101111;
				8'b111010: c <= 9'b1010011;
				8'b110110: c <= 9'b10101000;
				8'b1100100: c <= 9'b100001100;
				8'b1000000: c <= 9'b11111;
				8'b1110110: c <= 9'b10111100;
				8'b100101: c <= 9'b1001001;
				8'b101111: c <= 9'b101010101;
				8'b100110: c <= 9'b101111010;
				8'b1100011: c <= 9'b1101100;
				8'b1001000: c <= 9'b110001001;
				8'b111000: c <= 9'b10000001;
				8'b110001: c <= 9'b1010101;
				8'b1010111: c <= 9'b101010001;
				8'b1001110: c <= 9'b11001111;
				8'b1101010: c <= 9'b1000110;
				8'b1001001: c <= 9'b11100111;
				8'b1100000: c <= 9'b101011001;
				8'b110111: c <= 9'b100010110;
				8'b1011101: c <= 9'b111011001;
				8'b1011011: c <= 9'b100110110;
				8'b111001: c <= 9'b111000011;
				8'b1001010: c <= 9'b110100010;
				8'b110011: c <= 9'b1101010;
				8'b1101100: c <= 9'b110010001;
				8'b1110111: c <= 9'b1010000;
				8'b101011: c <= 9'b11;
				8'b1101011: c <= 9'b1101100;
				8'b111100: c <= 9'b11101101;
				8'b1000111: c <= 9'b1101010;
				8'b1011111: c <= 9'b11000011;
				8'b1110100: c <= 9'b110111110;
				8'b101101: c <= 9'b11000110;
				8'b1010011: c <= 9'b111101100;
				8'b1100001: c <= 9'b101101101;
				8'b110101: c <= 9'b111100011;
				8'b1000100: c <= 9'b100110;
				8'b1010001: c <= 9'b111001;
				8'b1010100: c <= 9'b110110110;
				8'b1100110: c <= 9'b111111111;
				8'b101010: c <= 9'b10100110;
				8'b1011110: c <= 9'b100001110;
				8'b1100111: c <= 9'b101010011;
				8'b1011010: c <= 9'b100101111;
				8'b1000010: c <= 9'b101110011;
				8'b111101: c <= 9'b110011;
				8'b110000: c <= 9'b110011;
				8'b111110: c <= 9'b101000;
				8'b1100010: c <= 9'b110000001;
				8'b1110000: c <= 9'b110001010;
				8'b1101001: c <= 9'b110101100;
				8'b1110011: c <= 9'b10011010;
				8'b1001100: c <= 9'b101000001;
				8'b100001: c <= 9'b11001111;
				8'b1000110: c <= 9'b10101010;
				8'b1110010: c <= 9'b11111100;
				8'b1010000: c <= 9'b100111111;
				8'b1111010: c <= 9'b100110110;
				8'b1010101: c <= 9'b100001110;
				8'b111011: c <= 9'b11101011;
				8'b1001101: c <= 9'b11000010;
				8'b111111: c <= 9'b1111111;
				8'b1101110: c <= 9'b10101;
				8'b1111011: c <= 9'b1101001;
				8'b1001011: c <= 9'b111000101;
				8'b1101111: c <= 9'b10010100;
				8'b1101000: c <= 9'b101001001;
				8'b101100: c <= 9'b110011000;
				8'b100100: c <= 9'b1001001;
				8'b1111000: c <= 9'b110110110;
				8'b1000101: c <= 9'b1001101;
				8'b1011001: c <= 9'b10101;
				8'b110100: c <= 9'b11111;
				8'b1111001: c <= 9'b1111111;
				8'b1110001: c <= 9'b111101111;
				8'b1001111: c <= 9'b101110101;
				8'b1100101: c <= 9'b10001001;
				8'b1111110: c <= 9'b101111110;
				8'b1111100: c <= 9'b1111011;
				8'b1010110: c <= 9'b10101011;
				8'b110010: c <= 9'b111000110;
				8'b1101101: c <= 9'b11101100;
				8'b100011: c <= 9'b100001101;
				8'b1110101: c <= 9'b11101100;
				8'b1111101: c <= 9'b1001;
				8'b101001: c <= 9'b100100011;
				8'b1010010: c <= 9'b110111000;
				8'b1011000: c <= 9'b101110010;
				8'b101110: c <= 9'b11000000;
				8'b1000001: c <= 9'b1011001;
				default: c <= 9'b0;
			endcase
			9'b1101010 : case(di)
				8'b1000011: c <= 9'b1100110;
				8'b101000: c <= 9'b100011001;
				8'b111010: c <= 9'b101010011;
				8'b110110: c <= 9'b11111001;
				8'b1100100: c <= 9'b101100;
				8'b1000000: c <= 9'b11000110;
				8'b1110110: c <= 9'b11010011;
				8'b100101: c <= 9'b1000100;
				8'b101111: c <= 9'b100000100;
				8'b100110: c <= 9'b100011101;
				8'b1100011: c <= 9'b11;
				8'b1001000: c <= 9'b110110100;
				8'b111000: c <= 9'b100111011;
				8'b110001: c <= 9'b110101101;
				8'b1010111: c <= 9'b110001011;
				8'b1001110: c <= 9'b110100011;
				8'b1101010: c <= 9'b1100;
				8'b1001001: c <= 9'b11011100;
				8'b1100000: c <= 9'b1000111;
				8'b110111: c <= 9'b101100110;
				8'b1011101: c <= 9'b100001001;
				8'b1011011: c <= 9'b11;
				8'b111001: c <= 9'b111111101;
				8'b1001010: c <= 9'b101100;
				8'b110011: c <= 9'b110101011;
				8'b1101100: c <= 9'b10100111;
				8'b1110111: c <= 9'b111100101;
				8'b101011: c <= 9'b11100000;
				8'b1101011: c <= 9'b100110011;
				8'b111100: c <= 9'b100101;
				8'b1000111: c <= 9'b100010010;
				8'b1011111: c <= 9'b11100;
				8'b1110100: c <= 9'b110101111;
				8'b101101: c <= 9'b111001010;
				8'b1010011: c <= 9'b1100101;
				8'b1100001: c <= 9'b101000010;
				8'b110101: c <= 9'b100000000;
				8'b1000100: c <= 9'b10010000;
				8'b1010001: c <= 9'b10011100;
				8'b1010100: c <= 9'b111111010;
				8'b1100110: c <= 9'b101101000;
				8'b101010: c <= 9'b11011;
				8'b1011110: c <= 9'b110110;
				8'b1100111: c <= 9'b100111000;
				8'b1011010: c <= 9'b111;
				8'b1000010: c <= 9'b111001;
				8'b111101: c <= 9'b1010010;
				8'b110000: c <= 9'b100101010;
				8'b111110: c <= 9'b110001001;
				8'b1100010: c <= 9'b1001010;
				8'b1110000: c <= 9'b100001111;
				8'b1101001: c <= 9'b11100011;
				8'b1110011: c <= 9'b1101110;
				8'b1001100: c <= 9'b1100100;
				8'b100001: c <= 9'b110110011;
				8'b1000110: c <= 9'b110111;
				8'b1110010: c <= 9'b10100101;
				8'b1010000: c <= 9'b100010101;
				8'b1111010: c <= 9'b11011100;
				8'b1010101: c <= 9'b101001001;
				8'b111011: c <= 9'b111001110;
				8'b1001101: c <= 9'b101010001;
				8'b111111: c <= 9'b110101111;
				8'b1101110: c <= 9'b1000101;
				8'b1111011: c <= 9'b10000101;
				8'b1001011: c <= 9'b1110011;
				8'b1101111: c <= 9'b100100111;
				8'b1101000: c <= 9'b111011100;
				8'b101100: c <= 9'b100111001;
				8'b100100: c <= 9'b110110100;
				8'b1111000: c <= 9'b110011101;
				8'b1000101: c <= 9'b10110101;
				8'b1011001: c <= 9'b1010010;
				8'b110100: c <= 9'b110100010;
				8'b1111001: c <= 9'b101000101;
				8'b1110001: c <= 9'b10111111;
				8'b1001111: c <= 9'b10011000;
				8'b1100101: c <= 9'b111001110;
				8'b1111110: c <= 9'b111011111;
				8'b1111100: c <= 9'b11011110;
				8'b1010110: c <= 9'b11100101;
				8'b110010: c <= 9'b101001;
				8'b1101101: c <= 9'b101001001;
				8'b100011: c <= 9'b111111011;
				8'b1110101: c <= 9'b10111011;
				8'b1111101: c <= 9'b100110111;
				8'b101001: c <= 9'b10010000;
				8'b1010010: c <= 9'b1101111;
				8'b1011000: c <= 9'b101001110;
				8'b101110: c <= 9'b1011110;
				8'b1000001: c <= 9'b101100;
				default: c <= 9'b0;
			endcase
			9'b1011010 : case(di)
				8'b1000011: c <= 9'b110011110;
				8'b101000: c <= 9'b101110010;
				8'b111010: c <= 9'b110010111;
				8'b110110: c <= 9'b10001110;
				8'b1100100: c <= 9'b11101;
				8'b1000000: c <= 9'b10110101;
				8'b1110110: c <= 9'b110001000;
				8'b100101: c <= 9'b10110111;
				8'b101111: c <= 9'b111101100;
				8'b100110: c <= 9'b101110101;
				8'b1100011: c <= 9'b100110110;
				8'b1001000: c <= 9'b101110010;
				8'b111000: c <= 9'b100100000;
				8'b110001: c <= 9'b110011000;
				8'b1010111: c <= 9'b1000110;
				8'b1001110: c <= 9'b100111001;
				8'b1101010: c <= 9'b101011110;
				8'b1001001: c <= 9'b100001001;
				8'b1100000: c <= 9'b1110111;
				8'b110111: c <= 9'b11111011;
				8'b1011101: c <= 9'b11101111;
				8'b1011011: c <= 9'b10001000;
				8'b111001: c <= 9'b100010101;
				8'b1001010: c <= 9'b10000101;
				8'b110011: c <= 9'b1001101;
				8'b1101100: c <= 9'b111010001;
				8'b1110111: c <= 9'b110100101;
				8'b101011: c <= 9'b11111110;
				8'b1101011: c <= 9'b110010;
				8'b111100: c <= 9'b110110100;
				8'b1000111: c <= 9'b10001111;
				8'b1011111: c <= 9'b11001111;
				8'b1110100: c <= 9'b101111110;
				8'b101101: c <= 9'b110111001;
				8'b1010011: c <= 9'b11000110;
				8'b1100001: c <= 9'b1011111;
				8'b110101: c <= 9'b10000010;
				8'b1000100: c <= 9'b111001110;
				8'b1010001: c <= 9'b101101000;
				8'b1010100: c <= 9'b110110011;
				8'b1100110: c <= 9'b111101110;
				8'b101010: c <= 9'b101000110;
				8'b1011110: c <= 9'b110101011;
				8'b1100111: c <= 9'b1000000;
				8'b1011010: c <= 9'b11001011;
				8'b1000010: c <= 9'b111110101;
				8'b111101: c <= 9'b100100001;
				8'b110000: c <= 9'b10011011;
				8'b111110: c <= 9'b111111111;
				8'b1100010: c <= 9'b11111011;
				8'b1110000: c <= 9'b100010001;
				8'b1101001: c <= 9'b11110110;
				8'b1110011: c <= 9'b11001000;
				8'b1001100: c <= 9'b11010010;
				8'b100001: c <= 9'b11100001;
				8'b1000110: c <= 9'b101111111;
				8'b1110010: c <= 9'b111111111;
				8'b1010000: c <= 9'b110011;
				8'b1111010: c <= 9'b101010001;
				8'b1010101: c <= 9'b11100111;
				8'b111011: c <= 9'b101100110;
				8'b1001101: c <= 9'b10111010;
				8'b111111: c <= 9'b100101000;
				8'b1101110: c <= 9'b101110011;
				8'b1111011: c <= 9'b100111000;
				8'b1001011: c <= 9'b10110101;
				8'b1101111: c <= 9'b11100;
				8'b1101000: c <= 9'b10111001;
				8'b101100: c <= 9'b100010110;
				8'b100100: c <= 9'b100000011;
				8'b1111000: c <= 9'b100110010;
				8'b1000101: c <= 9'b110001101;
				8'b1011001: c <= 9'b110010010;
				8'b110100: c <= 9'b110111110;
				8'b1111001: c <= 9'b1011001;
				8'b1110001: c <= 9'b10110010;
				8'b1001111: c <= 9'b101110111;
				8'b1100101: c <= 9'b110111110;
				8'b1111110: c <= 9'b101000001;
				8'b1111100: c <= 9'b10100100;
				8'b1010110: c <= 9'b11010101;
				8'b110010: c <= 9'b111100101;
				8'b1101101: c <= 9'b111100001;
				8'b100011: c <= 9'b11100111;
				8'b1110101: c <= 9'b11001;
				8'b1111101: c <= 9'b10001001;
				8'b101001: c <= 9'b110110100;
				8'b1010010: c <= 9'b100001010;
				8'b1011000: c <= 9'b1110000;
				8'b101110: c <= 9'b1000;
				8'b1000001: c <= 9'b110100101;
				default: c <= 9'b0;
			endcase
			9'b11110111 : case(di)
				8'b1000011: c <= 9'b111110000;
				8'b101000: c <= 9'b100011;
				8'b111010: c <= 9'b110111;
				8'b110110: c <= 9'b1010111;
				8'b1100100: c <= 9'b100010110;
				8'b1000000: c <= 9'b111110001;
				8'b1110110: c <= 9'b1011;
				8'b100101: c <= 9'b1110011;
				8'b101111: c <= 9'b11;
				8'b100110: c <= 9'b110100111;
				8'b1100011: c <= 9'b11111;
				8'b1001000: c <= 9'b100011100;
				8'b111000: c <= 9'b1111001;
				8'b110001: c <= 9'b110010001;
				8'b1010111: c <= 9'b10111010;
				8'b1001110: c <= 9'b111101100;
				8'b1101010: c <= 9'b10111101;
				8'b1001001: c <= 9'b1111101;
				8'b1100000: c <= 9'b1001010;
				8'b110111: c <= 9'b111011101;
				8'b1011101: c <= 9'b1111010;
				8'b1011011: c <= 9'b10111001;
				8'b111001: c <= 9'b11101000;
				8'b1001010: c <= 9'b1111100;
				8'b110011: c <= 9'b101001111;
				8'b1101100: c <= 9'b101010011;
				8'b1110111: c <= 9'b100011111;
				8'b101011: c <= 9'b1000010;
				8'b1101011: c <= 9'b11010010;
				8'b111100: c <= 9'b110;
				8'b1000111: c <= 9'b101000111;
				8'b1011111: c <= 9'b11100100;
				8'b1110100: c <= 9'b100010101;
				8'b101101: c <= 9'b110001010;
				8'b1010011: c <= 9'b100100011;
				8'b1100001: c <= 9'b110;
				8'b110101: c <= 9'b11111;
				8'b1000100: c <= 9'b101101111;
				8'b1010001: c <= 9'b110000111;
				8'b1010100: c <= 9'b101010000;
				8'b1100110: c <= 9'b1110011;
				8'b101010: c <= 9'b110111110;
				8'b1011110: c <= 9'b111000000;
				8'b1100111: c <= 9'b10100;
				8'b1011010: c <= 9'b111;
				8'b1000010: c <= 9'b1100;
				8'b111101: c <= 9'b111000110;
				8'b110000: c <= 9'b11010100;
				8'b111110: c <= 9'b1111111;
				8'b1100010: c <= 9'b111100111;
				8'b1110000: c <= 9'b10111101;
				8'b1101001: c <= 9'b110101101;
				8'b1110011: c <= 9'b101001001;
				8'b1001100: c <= 9'b110001000;
				8'b100001: c <= 9'b1111110;
				8'b1000110: c <= 9'b1101010;
				8'b1110010: c <= 9'b1110010;
				8'b1010000: c <= 9'b110001101;
				8'b1111010: c <= 9'b101100000;
				8'b1010101: c <= 9'b11011001;
				8'b111011: c <= 9'b10011100;
				8'b1001101: c <= 9'b1111001;
				8'b111111: c <= 9'b111010110;
				8'b1101110: c <= 9'b11011100;
				8'b1111011: c <= 9'b1011111;
				8'b1001011: c <= 9'b10100;
				8'b1101111: c <= 9'b11111010;
				8'b1101000: c <= 9'b10001101;
				8'b101100: c <= 9'b101000101;
				8'b100100: c <= 9'b110010;
				8'b1111000: c <= 9'b110000010;
				8'b1000101: c <= 9'b111011010;
				8'b1011001: c <= 9'b1000000;
				8'b110100: c <= 9'b10110100;
				8'b1111001: c <= 9'b110010110;
				8'b1110001: c <= 9'b11011101;
				8'b1001111: c <= 9'b111000011;
				8'b1100101: c <= 9'b1101101;
				8'b1111110: c <= 9'b1110;
				8'b1111100: c <= 9'b101101000;
				8'b1010110: c <= 9'b100001001;
				8'b110010: c <= 9'b101010010;
				8'b1101101: c <= 9'b10111001;
				8'b100011: c <= 9'b11100100;
				8'b1110101: c <= 9'b100100010;
				8'b1111101: c <= 9'b10011100;
				8'b101001: c <= 9'b11110;
				8'b1010010: c <= 9'b10;
				8'b1011000: c <= 9'b100001111;
				8'b101110: c <= 9'b11011001;
				8'b1000001: c <= 9'b10011010;
				default: c <= 9'b0;
			endcase
			9'b101101001 : case(di)
				8'b1000011: c <= 9'b100100001;
				8'b101000: c <= 9'b10010011;
				8'b111010: c <= 9'b100011101;
				8'b110110: c <= 9'b11110000;
				8'b1100100: c <= 9'b10101000;
				8'b1000000: c <= 9'b10100000;
				8'b1110110: c <= 9'b1100;
				8'b100101: c <= 9'b1001111;
				8'b101111: c <= 9'b101;
				8'b100110: c <= 9'b10011001;
				8'b1100011: c <= 9'b111010111;
				8'b1001000: c <= 9'b110010101;
				8'b111000: c <= 9'b101001;
				8'b110001: c <= 9'b110000111;
				8'b1010111: c <= 9'b100011011;
				8'b1001110: c <= 9'b10000101;
				8'b1101010: c <= 9'b10000101;
				8'b1001001: c <= 9'b101001100;
				8'b1100000: c <= 9'b1001;
				8'b110111: c <= 9'b10011010;
				8'b1011101: c <= 9'b110111001;
				8'b1011011: c <= 9'b111100110;
				8'b111001: c <= 9'b1101000;
				8'b1001010: c <= 9'b101111110;
				8'b110011: c <= 9'b11001;
				8'b1101100: c <= 9'b1000111;
				8'b1110111: c <= 9'b100000100;
				8'b101011: c <= 9'b101011111;
				8'b1101011: c <= 9'b1111100;
				8'b111100: c <= 9'b110001010;
				8'b1000111: c <= 9'b10101101;
				8'b1011111: c <= 9'b110110101;
				8'b1110100: c <= 9'b100010101;
				8'b101101: c <= 9'b110101011;
				8'b1010011: c <= 9'b100110111;
				8'b1100001: c <= 9'b100001100;
				8'b110101: c <= 9'b111100111;
				8'b1000100: c <= 9'b1010010;
				8'b1010001: c <= 9'b110110100;
				8'b1010100: c <= 9'b111100011;
				8'b1100110: c <= 9'b1010010;
				8'b101010: c <= 9'b11110100;
				8'b1011110: c <= 9'b11000110;
				8'b1100111: c <= 9'b11001;
				8'b1011010: c <= 9'b100011101;
				8'b1000010: c <= 9'b101001001;
				8'b111101: c <= 9'b101010001;
				8'b110000: c <= 9'b1111;
				8'b111110: c <= 9'b101001100;
				8'b1100010: c <= 9'b10001110;
				8'b1110000: c <= 9'b110000000;
				8'b1101001: c <= 9'b11011;
				8'b1110011: c <= 9'b101010110;
				8'b1001100: c <= 9'b111100;
				8'b100001: c <= 9'b101000100;
				8'b1000110: c <= 9'b100001111;
				8'b1110010: c <= 9'b111001111;
				8'b1010000: c <= 9'b110000110;
				8'b1111010: c <= 9'b11010011;
				8'b1010101: c <= 9'b10011100;
				8'b111011: c <= 9'b10011100;
				8'b1001101: c <= 9'b11100011;
				8'b111111: c <= 9'b100001110;
				8'b1101110: c <= 9'b1011011;
				8'b1111011: c <= 9'b111001100;
				8'b1001011: c <= 9'b110001011;
				8'b1101111: c <= 9'b11011101;
				8'b1101000: c <= 9'b101101110;
				8'b101100: c <= 9'b11001;
				8'b100100: c <= 9'b100001101;
				8'b1111000: c <= 9'b11000;
				8'b1000101: c <= 9'b11000100;
				8'b1011001: c <= 9'b101100000;
				8'b110100: c <= 9'b100010011;
				8'b1111001: c <= 9'b10110011;
				8'b1110001: c <= 9'b11110101;
				8'b1001111: c <= 9'b1000100;
				8'b1100101: c <= 9'b101100000;
				8'b1111110: c <= 9'b1001010;
				8'b1111100: c <= 9'b111111010;
				8'b1010110: c <= 9'b100011010;
				8'b110010: c <= 9'b111010001;
				8'b1101101: c <= 9'b101010101;
				8'b100011: c <= 9'b111110011;
				8'b1110101: c <= 9'b101001000;
				8'b1111101: c <= 9'b1100101;
				8'b101001: c <= 9'b1110011;
				8'b1010010: c <= 9'b10111001;
				8'b1011000: c <= 9'b100000001;
				8'b101110: c <= 9'b101011;
				8'b1000001: c <= 9'b110101;
				default: c <= 9'b0;
			endcase
			9'b10000000 : case(di)
				8'b1000011: c <= 9'b11011011;
				8'b101000: c <= 9'b100010;
				8'b111010: c <= 9'b10010001;
				8'b110110: c <= 9'b10100101;
				8'b1100100: c <= 9'b10101;
				8'b1000000: c <= 9'b10010101;
				8'b1110110: c <= 9'b111101010;
				8'b100101: c <= 9'b110000;
				8'b101111: c <= 9'b1011001;
				8'b100110: c <= 9'b111011001;
				8'b1100011: c <= 9'b11011011;
				8'b1001000: c <= 9'b111110001;
				8'b111000: c <= 9'b111000111;
				8'b110001: c <= 9'b111101111;
				8'b1010111: c <= 9'b100;
				8'b1001110: c <= 9'b11001000;
				8'b1101010: c <= 9'b101100111;
				8'b1001001: c <= 9'b111010111;
				8'b1100000: c <= 9'b101011;
				8'b110111: c <= 9'b100000110;
				8'b1011101: c <= 9'b10110111;
				8'b1011011: c <= 9'b101000110;
				8'b111001: c <= 9'b110101;
				8'b1001010: c <= 9'b11000100;
				8'b110011: c <= 9'b11011101;
				8'b1101100: c <= 9'b101000111;
				8'b1110111: c <= 9'b100010000;
				8'b101011: c <= 9'b11011100;
				8'b1101011: c <= 9'b11011000;
				8'b111100: c <= 9'b110001110;
				8'b1000111: c <= 9'b1100100;
				8'b1011111: c <= 9'b11011010;
				8'b1110100: c <= 9'b101101000;
				8'b101101: c <= 9'b10000010;
				8'b1010011: c <= 9'b101011011;
				8'b1100001: c <= 9'b11100110;
				8'b110101: c <= 9'b101010000;
				8'b1000100: c <= 9'b110111001;
				8'b1010001: c <= 9'b100100011;
				8'b1010100: c <= 9'b110101011;
				8'b1100110: c <= 9'b10100011;
				8'b101010: c <= 9'b10000111;
				8'b1011110: c <= 9'b11010010;
				8'b1100111: c <= 9'b11101;
				8'b1011010: c <= 9'b10010100;
				8'b1000010: c <= 9'b110001000;
				8'b111101: c <= 9'b1001101;
				8'b110000: c <= 9'b10001001;
				8'b111110: c <= 9'b10110110;
				8'b1100010: c <= 9'b111110001;
				8'b1110000: c <= 9'b10000111;
				8'b1101001: c <= 9'b111001101;
				8'b1110011: c <= 9'b110001;
				8'b1001100: c <= 9'b1111110;
				8'b100001: c <= 9'b10110101;
				8'b1000110: c <= 9'b11000000;
				8'b1110010: c <= 9'b101110010;
				8'b1010000: c <= 9'b11010001;
				8'b1111010: c <= 9'b111011100;
				8'b1010101: c <= 9'b1101100;
				8'b111011: c <= 9'b1000010;
				8'b1001101: c <= 9'b10000111;
				8'b111111: c <= 9'b1001001;
				8'b1101110: c <= 9'b11101011;
				8'b1111011: c <= 9'b101100111;
				8'b1001011: c <= 9'b110111;
				8'b1101111: c <= 9'b10110111;
				8'b1101000: c <= 9'b100101111;
				8'b101100: c <= 9'b110001011;
				8'b100100: c <= 9'b111100101;
				8'b1111000: c <= 9'b110101001;
				8'b1000101: c <= 9'b11010;
				8'b1011001: c <= 9'b100000111;
				8'b110100: c <= 9'b101110111;
				8'b1111001: c <= 9'b111010100;
				8'b1110001: c <= 9'b111101101;
				8'b1001111: c <= 9'b1100000;
				8'b1100101: c <= 9'b101001100;
				8'b1111110: c <= 9'b100010110;
				8'b1111100: c <= 9'b11101101;
				8'b1010110: c <= 9'b1100010;
				8'b110010: c <= 9'b10100000;
				8'b1101101: c <= 9'b10000111;
				8'b100011: c <= 9'b111010001;
				8'b1110101: c <= 9'b110000010;
				8'b1111101: c <= 9'b100011000;
				8'b101001: c <= 9'b100111001;
				8'b1010010: c <= 9'b110100110;
				8'b1011000: c <= 9'b111111011;
				8'b101110: c <= 9'b100111110;
				8'b1000001: c <= 9'b10001111;
				default: c <= 9'b0;
			endcase
			9'b101001110 : case(di)
				8'b1000011: c <= 9'b110110000;
				8'b101000: c <= 9'b100010101;
				8'b111010: c <= 9'b10010001;
				8'b110110: c <= 9'b101110001;
				8'b1100100: c <= 9'b11100101;
				8'b1000000: c <= 9'b101010011;
				8'b1110110: c <= 9'b101101011;
				8'b100101: c <= 9'b1000;
				8'b101111: c <= 9'b11011;
				8'b100110: c <= 9'b10101010;
				8'b1100011: c <= 9'b100000110;
				8'b1001000: c <= 9'b1;
				8'b111000: c <= 9'b11101101;
				8'b110001: c <= 9'b10111101;
				8'b1010111: c <= 9'b10110001;
				8'b1001110: c <= 9'b111011011;
				8'b1101010: c <= 9'b111001101;
				8'b1001001: c <= 9'b1000001;
				8'b1100000: c <= 9'b111010100;
				8'b110111: c <= 9'b10010011;
				8'b1011101: c <= 9'b1011111;
				8'b1011011: c <= 9'b110000011;
				8'b111001: c <= 9'b110100;
				8'b1001010: c <= 9'b11000;
				8'b110011: c <= 9'b10011101;
				8'b1101100: c <= 9'b111010000;
				8'b1110111: c <= 9'b11010100;
				8'b101011: c <= 9'b100101111;
				8'b1101011: c <= 9'b111111000;
				8'b111100: c <= 9'b101011001;
				8'b1000111: c <= 9'b1100101;
				8'b1011111: c <= 9'b100101101;
				8'b1110100: c <= 9'b110111010;
				8'b101101: c <= 9'b1101100;
				8'b1010011: c <= 9'b1101;
				8'b1100001: c <= 9'b10000001;
				8'b110101: c <= 9'b11011011;
				8'b1000100: c <= 9'b111001111;
				8'b1010001: c <= 9'b10110001;
				8'b1010100: c <= 9'b111100000;
				8'b1100110: c <= 9'b110001111;
				8'b101010: c <= 9'b110011101;
				8'b1011110: c <= 9'b1101111;
				8'b1100111: c <= 9'b101111010;
				8'b1011010: c <= 9'b1101001;
				8'b1000010: c <= 9'b110001111;
				8'b111101: c <= 9'b11110100;
				8'b110000: c <= 9'b1100001;
				8'b111110: c <= 9'b10100101;
				8'b1100010: c <= 9'b11110;
				8'b1110000: c <= 9'b110111000;
				8'b1101001: c <= 9'b1000001;
				8'b1110011: c <= 9'b1011110;
				8'b1001100: c <= 9'b101001001;
				8'b100001: c <= 9'b111010;
				8'b1000110: c <= 9'b111111;
				8'b1110010: c <= 9'b111100100;
				8'b1010000: c <= 9'b101011001;
				8'b1111010: c <= 9'b11100000;
				8'b1010101: c <= 9'b101011010;
				8'b111011: c <= 9'b111101;
				8'b1001101: c <= 9'b100011001;
				8'b111111: c <= 9'b110111010;
				8'b1101110: c <= 9'b110111000;
				8'b1111011: c <= 9'b110101100;
				8'b1001011: c <= 9'b101011111;
				8'b1101111: c <= 9'b101110010;
				8'b1101000: c <= 9'b101111111;
				8'b101100: c <= 9'b110011111;
				8'b100100: c <= 9'b101110111;
				8'b1111000: c <= 9'b11111110;
				8'b1000101: c <= 9'b11111100;
				8'b1011001: c <= 9'b11111000;
				8'b110100: c <= 9'b10111111;
				8'b1111001: c <= 9'b11010111;
				8'b1110001: c <= 9'b100001011;
				8'b1001111: c <= 9'b10000000;
				8'b1100101: c <= 9'b111011001;
				8'b1111110: c <= 9'b110000111;
				8'b1111100: c <= 9'b10001010;
				8'b1010110: c <= 9'b11001111;
				8'b110010: c <= 9'b111100111;
				8'b1101101: c <= 9'b11000100;
				8'b100011: c <= 9'b111010111;
				8'b1110101: c <= 9'b101110010;
				8'b1111101: c <= 9'b10011100;
				8'b101001: c <= 9'b101101100;
				8'b1010010: c <= 9'b10001001;
				8'b1011000: c <= 9'b11101;
				8'b101110: c <= 9'b100100101;
				8'b1000001: c <= 9'b110001111;
				default: c <= 9'b0;
			endcase
			9'b110011 : case(di)
				8'b1000011: c <= 9'b11010010;
				8'b101000: c <= 9'b111010100;
				8'b111010: c <= 9'b101010011;
				8'b110110: c <= 9'b10000001;
				8'b1100100: c <= 9'b11011000;
				8'b1000000: c <= 9'b10110010;
				8'b1110110: c <= 9'b100010110;
				8'b100101: c <= 9'b1010010;
				8'b101111: c <= 9'b111000;
				8'b100110: c <= 9'b100111111;
				8'b1100011: c <= 9'b110000011;
				8'b1001000: c <= 9'b100011;
				8'b111000: c <= 9'b100011;
				8'b110001: c <= 9'b1000110;
				8'b1010111: c <= 9'b11110010;
				8'b1001110: c <= 9'b111010;
				8'b1101010: c <= 9'b111110001;
				8'b1001001: c <= 9'b1101000;
				8'b1100000: c <= 9'b101110011;
				8'b110111: c <= 9'b111101100;
				8'b1011101: c <= 9'b111101100;
				8'b1011011: c <= 9'b110010011;
				8'b111001: c <= 9'b11110101;
				8'b1001010: c <= 9'b10101101;
				8'b110011: c <= 9'b100010100;
				8'b1101100: c <= 9'b1101;
				8'b1110111: c <= 9'b101101010;
				8'b101011: c <= 9'b110110101;
				8'b1101011: c <= 9'b10100111;
				8'b111100: c <= 9'b111000111;
				8'b1000111: c <= 9'b10100101;
				8'b1011111: c <= 9'b101111010;
				8'b1110100: c <= 9'b1101;
				8'b101101: c <= 9'b10101111;
				8'b1010011: c <= 9'b110010011;
				8'b1100001: c <= 9'b1001111;
				8'b110101: c <= 9'b10000011;
				8'b1000100: c <= 9'b100000011;
				8'b1010001: c <= 9'b10001101;
				8'b1010100: c <= 9'b111001011;
				8'b1100110: c <= 9'b111001000;
				8'b101010: c <= 9'b101001100;
				8'b1011110: c <= 9'b111001000;
				8'b1100111: c <= 9'b1111110;
				8'b1011010: c <= 9'b101001;
				8'b1000010: c <= 9'b111100;
				8'b111101: c <= 9'b100101111;
				8'b110000: c <= 9'b110010010;
				8'b111110: c <= 9'b101010011;
				8'b1100010: c <= 9'b101010011;
				8'b1110000: c <= 9'b101000011;
				8'b1101001: c <= 9'b101100;
				8'b1110011: c <= 9'b111000011;
				8'b1001100: c <= 9'b101010001;
				8'b100001: c <= 9'b101110;
				8'b1000110: c <= 9'b11011101;
				8'b1110010: c <= 9'b1110001;
				8'b1010000: c <= 9'b10101000;
				8'b1111010: c <= 9'b100010111;
				8'b1010101: c <= 9'b11110111;
				8'b111011: c <= 9'b111111101;
				8'b1001101: c <= 9'b100000110;
				8'b111111: c <= 9'b100100;
				8'b1101110: c <= 9'b111011011;
				8'b1111011: c <= 9'b11101000;
				8'b1001011: c <= 9'b110100000;
				8'b1101111: c <= 9'b111000100;
				8'b1101000: c <= 9'b10111011;
				8'b101100: c <= 9'b111101110;
				8'b100100: c <= 9'b10010;
				8'b1111000: c <= 9'b10111111;
				8'b1000101: c <= 9'b111110000;
				8'b1011001: c <= 9'b110010100;
				8'b110100: c <= 9'b1011010;
				8'b1111001: c <= 9'b111100001;
				8'b1110001: c <= 9'b11001101;
				8'b1001111: c <= 9'b111101101;
				8'b1100101: c <= 9'b10100;
				8'b1111110: c <= 9'b10001100;
				8'b1111100: c <= 9'b110100100;
				8'b1010110: c <= 9'b101110000;
				8'b110010: c <= 9'b10110100;
				8'b1101101: c <= 9'b111001010;
				8'b100011: c <= 9'b10111010;
				8'b1110101: c <= 9'b11010011;
				8'b1111101: c <= 9'b10110001;
				8'b101001: c <= 9'b11101;
				8'b1010010: c <= 9'b111101010;
				8'b1011000: c <= 9'b110000110;
				8'b101110: c <= 9'b100111101;
				8'b1000001: c <= 9'b110011100;
				default: c <= 9'b0;
			endcase
			9'b111010001 : case(di)
				8'b1000011: c <= 9'b1010001;
				8'b101000: c <= 9'b11001010;
				8'b111010: c <= 9'b11001001;
				8'b110110: c <= 9'b1000011;
				8'b1100100: c <= 9'b111101111;
				8'b1000000: c <= 9'b101111110;
				8'b1110110: c <= 9'b1110010;
				8'b100101: c <= 9'b11110001;
				8'b101111: c <= 9'b1111011;
				8'b100110: c <= 9'b1100110;
				8'b1100011: c <= 9'b100010111;
				8'b1001000: c <= 9'b1110100;
				8'b111000: c <= 9'b11101001;
				8'b110001: c <= 9'b11110001;
				8'b1010111: c <= 9'b11010100;
				8'b1001110: c <= 9'b111001000;
				8'b1101010: c <= 9'b1101000;
				8'b1001001: c <= 9'b101101101;
				8'b1100000: c <= 9'b100000111;
				8'b110111: c <= 9'b111011;
				8'b1011101: c <= 9'b110101001;
				8'b1011011: c <= 9'b11010100;
				8'b111001: c <= 9'b10000;
				8'b1001010: c <= 9'b10010;
				8'b110011: c <= 9'b110011;
				8'b1101100: c <= 9'b11101011;
				8'b1110111: c <= 9'b10101;
				8'b101011: c <= 9'b10111;
				8'b1101011: c <= 9'b111000111;
				8'b111100: c <= 9'b11010111;
				8'b1000111: c <= 9'b10110111;
				8'b1011111: c <= 9'b11011100;
				8'b1110100: c <= 9'b100100000;
				8'b101101: c <= 9'b110010001;
				8'b1010011: c <= 9'b1011110;
				8'b1100001: c <= 9'b10011100;
				8'b110101: c <= 9'b10111100;
				8'b1000100: c <= 9'b110011011;
				8'b1010001: c <= 9'b110011;
				8'b1010100: c <= 9'b1110011;
				8'b1100110: c <= 9'b100000011;
				8'b101010: c <= 9'b110110111;
				8'b1011110: c <= 9'b111100000;
				8'b1100111: c <= 9'b10101001;
				8'b1011010: c <= 9'b10000110;
				8'b1000010: c <= 9'b1101111;
				8'b111101: c <= 9'b11000;
				8'b110000: c <= 9'b10001010;
				8'b111110: c <= 9'b1111001;
				8'b1100010: c <= 9'b110110;
				8'b1110000: c <= 9'b110100000;
				8'b1101001: c <= 9'b111011111;
				8'b1110011: c <= 9'b111011010;
				8'b1001100: c <= 9'b100110;
				8'b100001: c <= 9'b11111000;
				8'b1000110: c <= 9'b110000010;
				8'b1110010: c <= 9'b11110000;
				8'b1010000: c <= 9'b1110011;
				8'b1111010: c <= 9'b100110101;
				8'b1010101: c <= 9'b1010010;
				8'b111011: c <= 9'b110110111;
				8'b1001101: c <= 9'b101101111;
				8'b111111: c <= 9'b11101001;
				8'b1101110: c <= 9'b101000010;
				8'b1111011: c <= 9'b110011;
				8'b1001011: c <= 9'b101010010;
				8'b1101111: c <= 9'b101011010;
				8'b1101000: c <= 9'b101000100;
				8'b101100: c <= 9'b11110110;
				8'b100100: c <= 9'b1111110;
				8'b1111000: c <= 9'b110001000;
				8'b1000101: c <= 9'b110011011;
				8'b1011001: c <= 9'b100000110;
				8'b110100: c <= 9'b10010000;
				8'b1111001: c <= 9'b11110110;
				8'b1110001: c <= 9'b10011000;
				8'b1001111: c <= 9'b100110100;
				8'b1100101: c <= 9'b10001101;
				8'b1111110: c <= 9'b1110011;
				8'b1111100: c <= 9'b111101001;
				8'b1010110: c <= 9'b11000110;
				8'b110010: c <= 9'b10110011;
				8'b1101101: c <= 9'b100011011;
				8'b100011: c <= 9'b111111011;
				8'b1110101: c <= 9'b100100001;
				8'b1111101: c <= 9'b111100010;
				8'b101001: c <= 9'b111011111;
				8'b1010010: c <= 9'b10011010;
				8'b1011000: c <= 9'b110110011;
				8'b101110: c <= 9'b11;
				8'b1000001: c <= 9'b101010000;
				default: c <= 9'b0;
			endcase
			9'b1000011 : case(di)
				8'b1000011: c <= 9'b110000110;
				8'b101000: c <= 9'b10110110;
				8'b111010: c <= 9'b101011111;
				8'b110110: c <= 9'b101000011;
				8'b1100100: c <= 9'b10100100;
				8'b1000000: c <= 9'b100010100;
				8'b1110110: c <= 9'b101100001;
				8'b100101: c <= 9'b110010110;
				8'b101111: c <= 9'b1101100;
				8'b100110: c <= 9'b10001110;
				8'b1100011: c <= 9'b10111101;
				8'b1001000: c <= 9'b10010001;
				8'b111000: c <= 9'b1100011;
				8'b110001: c <= 9'b101110100;
				8'b1010111: c <= 9'b101011;
				8'b1001110: c <= 9'b10000;
				8'b1101010: c <= 9'b1110011;
				8'b1001001: c <= 9'b1110011;
				8'b1100000: c <= 9'b111011101;
				8'b110111: c <= 9'b1110010;
				8'b1011101: c <= 9'b101110101;
				8'b1011011: c <= 9'b111101110;
				8'b111001: c <= 9'b111010100;
				8'b1001010: c <= 9'b110111110;
				8'b110011: c <= 9'b10001010;
				8'b1101100: c <= 9'b10110;
				8'b1110111: c <= 9'b1000111;
				8'b101011: c <= 9'b11001;
				8'b1101011: c <= 9'b110111001;
				8'b111100: c <= 9'b1000111;
				8'b1000111: c <= 9'b101010110;
				8'b1011111: c <= 9'b111011111;
				8'b1110100: c <= 9'b110010010;
				8'b101101: c <= 9'b1001111;
				8'b1010011: c <= 9'b110101110;
				8'b1100001: c <= 9'b1;
				8'b110101: c <= 9'b100111010;
				8'b1000100: c <= 9'b10101001;
				8'b1010001: c <= 9'b101010;
				8'b1010100: c <= 9'b100110011;
				8'b1100110: c <= 9'b111011010;
				8'b101010: c <= 9'b101011000;
				8'b1011110: c <= 9'b100101111;
				8'b1100111: c <= 9'b10110;
				8'b1011010: c <= 9'b111000000;
				8'b1000010: c <= 9'b100000111;
				8'b111101: c <= 9'b10001100;
				8'b110000: c <= 9'b1110100;
				8'b111110: c <= 9'b11110111;
				8'b1100010: c <= 9'b101010000;
				8'b1110000: c <= 9'b100110100;
				8'b1101001: c <= 9'b10001011;
				8'b1110011: c <= 9'b1011010;
				8'b1001100: c <= 9'b101110000;
				8'b100001: c <= 9'b100111111;
				8'b1000110: c <= 9'b110110101;
				8'b1110010: c <= 9'b101001100;
				8'b1010000: c <= 9'b101010100;
				8'b1111010: c <= 9'b111011101;
				8'b1010101: c <= 9'b110;
				8'b111011: c <= 9'b11010000;
				8'b1001101: c <= 9'b101010000;
				8'b111111: c <= 9'b10110010;
				8'b1101110: c <= 9'b101011010;
				8'b1111011: c <= 9'b111111110;
				8'b1001011: c <= 9'b10100010;
				8'b1101111: c <= 9'b11010100;
				8'b1101000: c <= 9'b110001;
				8'b101100: c <= 9'b101010000;
				8'b100100: c <= 9'b111110000;
				8'b1111000: c <= 9'b1111010;
				8'b1000101: c <= 9'b110011101;
				8'b1011001: c <= 9'b111010;
				8'b110100: c <= 9'b101100011;
				8'b1111001: c <= 9'b10;
				8'b1110001: c <= 9'b110111110;
				8'b1001111: c <= 9'b111001011;
				8'b1100101: c <= 9'b10111101;
				8'b1111110: c <= 9'b11100111;
				8'b1111100: c <= 9'b11011100;
				8'b1010110: c <= 9'b1101110;
				8'b110010: c <= 9'b10011000;
				8'b1101101: c <= 9'b10;
				8'b100011: c <= 9'b111001001;
				8'b1110101: c <= 9'b1010111;
				8'b1111101: c <= 9'b110001001;
				8'b101001: c <= 9'b11010100;
				8'b1010010: c <= 9'b100101001;
				8'b1011000: c <= 9'b100110100;
				8'b101110: c <= 9'b1100111;
				8'b1000001: c <= 9'b110100011;
				default: c <= 9'b0;
			endcase
			9'b111111010 : case(di)
				8'b1000011: c <= 9'b1101111;
				8'b101000: c <= 9'b1010010;
				8'b111010: c <= 9'b100011111;
				8'b110110: c <= 9'b11100011;
				8'b1100100: c <= 9'b100011010;
				8'b1000000: c <= 9'b110000001;
				8'b1110110: c <= 9'b11100001;
				8'b100101: c <= 9'b110100110;
				8'b101111: c <= 9'b100010110;
				8'b100110: c <= 9'b10100111;
				8'b1100011: c <= 9'b111100;
				8'b1001000: c <= 9'b11000100;
				8'b111000: c <= 9'b11101;
				8'b110001: c <= 9'b1001101;
				8'b1010111: c <= 9'b100010010;
				8'b1001110: c <= 9'b11111100;
				8'b1101010: c <= 9'b110100000;
				8'b1001001: c <= 9'b11100110;
				8'b1100000: c <= 9'b1000101;
				8'b110111: c <= 9'b101111110;
				8'b1011101: c <= 9'b101111111;
				8'b1011011: c <= 9'b1110;
				8'b111001: c <= 9'b11111010;
				8'b1001010: c <= 9'b111001000;
				8'b110011: c <= 9'b100101101;
				8'b1101100: c <= 9'b10001100;
				8'b1110111: c <= 9'b1111011;
				8'b101011: c <= 9'b101011101;
				8'b1101011: c <= 9'b111010100;
				8'b111100: c <= 9'b101110;
				8'b1000111: c <= 9'b101101011;
				8'b1011111: c <= 9'b111101110;
				8'b1110100: c <= 9'b101011010;
				8'b101101: c <= 9'b11010000;
				8'b1010011: c <= 9'b110101100;
				8'b1100001: c <= 9'b101001;
				8'b110101: c <= 9'b10011000;
				8'b1000100: c <= 9'b100000100;
				8'b1010001: c <= 9'b110011111;
				8'b1010100: c <= 9'b100110011;
				8'b1100110: c <= 9'b110010100;
				8'b101010: c <= 9'b101110;
				8'b1011110: c <= 9'b11100010;
				8'b1100111: c <= 9'b110011111;
				8'b1011010: c <= 9'b10000110;
				8'b1000010: c <= 9'b10110110;
				8'b111101: c <= 9'b101110111;
				8'b110000: c <= 9'b11100111;
				8'b111110: c <= 9'b10001110;
				8'b1100010: c <= 9'b11000;
				8'b1110000: c <= 9'b1110101;
				8'b1101001: c <= 9'b11010100;
				8'b1110011: c <= 9'b101111000;
				8'b1001100: c <= 9'b1100101;
				8'b100001: c <= 9'b101011000;
				8'b1000110: c <= 9'b1110111;
				8'b1110010: c <= 9'b111101111;
				8'b1010000: c <= 9'b101011111;
				8'b1111010: c <= 9'b10101101;
				8'b1010101: c <= 9'b110110110;
				8'b111011: c <= 9'b11011010;
				8'b1001101: c <= 9'b111110101;
				8'b111111: c <= 9'b10111101;
				8'b1101110: c <= 9'b1111010;
				8'b1111011: c <= 9'b1011000;
				8'b1001011: c <= 9'b111000110;
				8'b1101111: c <= 9'b101100110;
				8'b1101000: c <= 9'b100000111;
				8'b101100: c <= 9'b101000111;
				8'b100100: c <= 9'b11100111;
				8'b1111000: c <= 9'b101010;
				8'b1000101: c <= 9'b110110010;
				8'b1011001: c <= 9'b1100010;
				8'b110100: c <= 9'b110011110;
				8'b1111001: c <= 9'b111001100;
				8'b1110001: c <= 9'b11010001;
				8'b1001111: c <= 9'b1111111;
				8'b1100101: c <= 9'b1010001;
				8'b1111110: c <= 9'b1100010;
				8'b1111100: c <= 9'b100101111;
				8'b1010110: c <= 9'b101100111;
				8'b110010: c <= 9'b10100111;
				8'b1101101: c <= 9'b1000;
				8'b100011: c <= 9'b100001110;
				8'b1110101: c <= 9'b100110110;
				8'b1111101: c <= 9'b101000100;
				8'b101001: c <= 9'b110110000;
				8'b1010010: c <= 9'b1001100;
				8'b1011000: c <= 9'b10010101;
				8'b101110: c <= 9'b10100010;
				8'b1000001: c <= 9'b111001011;
				default: c <= 9'b0;
			endcase
			9'b100000110 : case(di)
				8'b1000011: c <= 9'b110011110;
				8'b101000: c <= 9'b10010110;
				8'b111010: c <= 9'b110000001;
				8'b110110: c <= 9'b101010010;
				8'b1100100: c <= 9'b101010010;
				8'b1000000: c <= 9'b11101100;
				8'b1110110: c <= 9'b110010110;
				8'b100101: c <= 9'b100000111;
				8'b101111: c <= 9'b11110;
				8'b100110: c <= 9'b1001110;
				8'b1100011: c <= 9'b10110111;
				8'b1001000: c <= 9'b101101011;
				8'b111000: c <= 9'b110101010;
				8'b110001: c <= 9'b110100110;
				8'b1010111: c <= 9'b10100110;
				8'b1001110: c <= 9'b11111100;
				8'b1101010: c <= 9'b10100100;
				8'b1001001: c <= 9'b11101000;
				8'b1100000: c <= 9'b10111101;
				8'b110111: c <= 9'b101000;
				8'b1011101: c <= 9'b10101100;
				8'b1011011: c <= 9'b11100111;
				8'b111001: c <= 9'b1001010;
				8'b1001010: c <= 9'b111010110;
				8'b110011: c <= 9'b111001;
				8'b1101100: c <= 9'b101110001;
				8'b1110111: c <= 9'b111000110;
				8'b101011: c <= 9'b101;
				8'b1101011: c <= 9'b110001010;
				8'b111100: c <= 9'b101001000;
				8'b1000111: c <= 9'b111010000;
				8'b1011111: c <= 9'b100110000;
				8'b1110100: c <= 9'b11010011;
				8'b101101: c <= 9'b1101010;
				8'b1010011: c <= 9'b100010110;
				8'b1100001: c <= 9'b10001101;
				8'b110101: c <= 9'b11111011;
				8'b1000100: c <= 9'b10101100;
				8'b1010001: c <= 9'b111011011;
				8'b1010100: c <= 9'b11010100;
				8'b1100110: c <= 9'b100111111;
				8'b101010: c <= 9'b111100000;
				8'b1011110: c <= 9'b11001110;
				8'b1100111: c <= 9'b100010010;
				8'b1011010: c <= 9'b11110101;
				8'b1000010: c <= 9'b110010111;
				8'b111101: c <= 9'b1110011;
				8'b110000: c <= 9'b110101011;
				8'b111110: c <= 9'b11111100;
				8'b1100010: c <= 9'b110010001;
				8'b1110000: c <= 9'b1101101;
				8'b1101001: c <= 9'b10001110;
				8'b1110011: c <= 9'b1111000;
				8'b1001100: c <= 9'b11100111;
				8'b100001: c <= 9'b101010101;
				8'b1000110: c <= 9'b1111;
				8'b1110010: c <= 9'b110001;
				8'b1010000: c <= 9'b10001001;
				8'b1111010: c <= 9'b100010101;
				8'b1010101: c <= 9'b110001111;
				8'b111011: c <= 9'b111101010;
				8'b1001101: c <= 9'b110101101;
				8'b111111: c <= 9'b100001001;
				8'b1101110: c <= 9'b11111010;
				8'b1111011: c <= 9'b10000111;
				8'b1001011: c <= 9'b100;
				8'b1101111: c <= 9'b100011111;
				8'b1101000: c <= 9'b100011100;
				8'b101100: c <= 9'b101101;
				8'b100100: c <= 9'b101101100;
				8'b1111000: c <= 9'b111001101;
				8'b1000101: c <= 9'b1011111;
				8'b1011001: c <= 9'b111110011;
				8'b110100: c <= 9'b101110010;
				8'b1111001: c <= 9'b10111;
				8'b1110001: c <= 9'b11100011;
				8'b1001111: c <= 9'b11010100;
				8'b1100101: c <= 9'b110110101;
				8'b1111110: c <= 9'b100010010;
				8'b1111100: c <= 9'b100111110;
				8'b1010110: c <= 9'b111011001;
				8'b110010: c <= 9'b1001;
				8'b1101101: c <= 9'b110001010;
				8'b100011: c <= 9'b11110110;
				8'b1110101: c <= 9'b110101111;
				8'b1111101: c <= 9'b110100011;
				8'b101001: c <= 9'b10110;
				8'b1010010: c <= 9'b111000111;
				8'b1011000: c <= 9'b110001000;
				8'b101110: c <= 9'b11001111;
				8'b1000001: c <= 9'b11000100;
				default: c <= 9'b0;
			endcase
			9'b100010000 : case(di)
				8'b1000011: c <= 9'b101101;
				8'b101000: c <= 9'b100000111;
				8'b111010: c <= 9'b1010111;
				8'b110110: c <= 9'b10100011;
				8'b1100100: c <= 9'b10001000;
				8'b1000000: c <= 9'b11100001;
				8'b1110110: c <= 9'b100000101;
				8'b100101: c <= 9'b110100111;
				8'b101111: c <= 9'b100101110;
				8'b100110: c <= 9'b110001100;
				8'b1100011: c <= 9'b1011100;
				8'b1001000: c <= 9'b111101;
				8'b111000: c <= 9'b10101001;
				8'b110001: c <= 9'b1111011;
				8'b1010111: c <= 9'b1010011;
				8'b1001110: c <= 9'b101100000;
				8'b1101010: c <= 9'b110011100;
				8'b1001001: c <= 9'b10010001;
				8'b1100000: c <= 9'b10111111;
				8'b110111: c <= 9'b1101101;
				8'b1011101: c <= 9'b101110;
				8'b1011011: c <= 9'b110011011;
				8'b111001: c <= 9'b1011100;
				8'b1001010: c <= 9'b11001011;
				8'b110011: c <= 9'b10101111;
				8'b1101100: c <= 9'b10010;
				8'b1110111: c <= 9'b10110;
				8'b101011: c <= 9'b110001101;
				8'b1101011: c <= 9'b1010010;
				8'b111100: c <= 9'b1000110;
				8'b1000111: c <= 9'b110001110;
				8'b1011111: c <= 9'b100;
				8'b1110100: c <= 9'b10101001;
				8'b101101: c <= 9'b1100001;
				8'b1010011: c <= 9'b101000010;
				8'b1100001: c <= 9'b100110111;
				8'b110101: c <= 9'b11100;
				8'b1000100: c <= 9'b110010110;
				8'b1010001: c <= 9'b101111111;
				8'b1010100: c <= 9'b1111100;
				8'b1100110: c <= 9'b110000111;
				8'b101010: c <= 9'b1010011;
				8'b1011110: c <= 9'b111110101;
				8'b1100111: c <= 9'b1000100;
				8'b1011010: c <= 9'b101001000;
				8'b1000010: c <= 9'b101000101;
				8'b111101: c <= 9'b100101101;
				8'b110000: c <= 9'b111000110;
				8'b111110: c <= 9'b11100000;
				8'b1100010: c <= 9'b111111010;
				8'b1110000: c <= 9'b101111001;
				8'b1101001: c <= 9'b100100101;
				8'b1110011: c <= 9'b111010010;
				8'b1001100: c <= 9'b11010010;
				8'b100001: c <= 9'b111111111;
				8'b1000110: c <= 9'b111001000;
				8'b1110010: c <= 9'b100000111;
				8'b1010000: c <= 9'b110000001;
				8'b1111010: c <= 9'b11000001;
				8'b1010101: c <= 9'b101001010;
				8'b111011: c <= 9'b1111110;
				8'b1001101: c <= 9'b110000010;
				8'b111111: c <= 9'b110110101;
				8'b1101110: c <= 9'b10101110;
				8'b1111011: c <= 9'b11101;
				8'b1001011: c <= 9'b100100001;
				8'b1101111: c <= 9'b100101010;
				8'b1101000: c <= 9'b10010111;
				8'b101100: c <= 9'b11001;
				8'b100100: c <= 9'b101101111;
				8'b1111000: c <= 9'b10100110;
				8'b1000101: c <= 9'b101001001;
				8'b1011001: c <= 9'b10;
				8'b110100: c <= 9'b100010;
				8'b1111001: c <= 9'b1011001;
				8'b1110001: c <= 9'b10;
				8'b1001111: c <= 9'b101011110;
				8'b1100101: c <= 9'b10111101;
				8'b1111110: c <= 9'b10110110;
				8'b1111100: c <= 9'b111111110;
				8'b1010110: c <= 9'b1010001;
				8'b110010: c <= 9'b10010001;
				8'b1101101: c <= 9'b110100100;
				8'b100011: c <= 9'b11101100;
				8'b1110101: c <= 9'b101000;
				8'b1111101: c <= 9'b110111110;
				8'b101001: c <= 9'b101100110;
				8'b1010010: c <= 9'b1100001;
				8'b1011000: c <= 9'b1101001;
				8'b101110: c <= 9'b10001001;
				8'b1000001: c <= 9'b110001001;
				default: c <= 9'b0;
			endcase
			9'b110011010 : case(di)
				8'b1000011: c <= 9'b100;
				8'b101000: c <= 9'b10000011;
				8'b111010: c <= 9'b110100111;
				8'b110110: c <= 9'b100101;
				8'b1100100: c <= 9'b111101010;
				8'b1000000: c <= 9'b101110110;
				8'b1110110: c <= 9'b101010100;
				8'b100101: c <= 9'b10100110;
				8'b101111: c <= 9'b111000111;
				8'b100110: c <= 9'b101001011;
				8'b1100011: c <= 9'b100100010;
				8'b1001000: c <= 9'b100111001;
				8'b111000: c <= 9'b11001;
				8'b110001: c <= 9'b10110010;
				8'b1010111: c <= 9'b100110100;
				8'b1001110: c <= 9'b11100100;
				8'b1101010: c <= 9'b101110001;
				8'b1001001: c <= 9'b101011;
				8'b1100000: c <= 9'b1011110;
				8'b110111: c <= 9'b111101101;
				8'b1011101: c <= 9'b11001011;
				8'b1011011: c <= 9'b10101111;
				8'b111001: c <= 9'b110111110;
				8'b1001010: c <= 9'b1110000;
				8'b110011: c <= 9'b111010110;
				8'b1101100: c <= 9'b100101101;
				8'b1110111: c <= 9'b101011111;
				8'b101011: c <= 9'b110111011;
				8'b1101011: c <= 9'b101111001;
				8'b111100: c <= 9'b111010110;
				8'b1000111: c <= 9'b11000110;
				8'b1011111: c <= 9'b111000101;
				8'b1110100: c <= 9'b110001011;
				8'b101101: c <= 9'b1101;
				8'b1010011: c <= 9'b100010001;
				8'b1100001: c <= 9'b101000101;
				8'b110101: c <= 9'b1111;
				8'b1000100: c <= 9'b101101001;
				8'b1010001: c <= 9'b10100000;
				8'b1010100: c <= 9'b11001100;
				8'b1100110: c <= 9'b100110101;
				8'b101010: c <= 9'b110101101;
				8'b1011110: c <= 9'b111000000;
				8'b1100111: c <= 9'b101100011;
				8'b1011010: c <= 9'b10001011;
				8'b1000010: c <= 9'b110101001;
				8'b111101: c <= 9'b110101;
				8'b110000: c <= 9'b101011111;
				8'b111110: c <= 9'b10001100;
				8'b1100010: c <= 9'b100000010;
				8'b1110000: c <= 9'b10110100;
				8'b1101001: c <= 9'b100111100;
				8'b1110011: c <= 9'b101111110;
				8'b1001100: c <= 9'b100111010;
				8'b100001: c <= 9'b110011001;
				8'b1000110: c <= 9'b101101001;
				8'b1110010: c <= 9'b110111010;
				8'b1010000: c <= 9'b100001010;
				8'b1111010: c <= 9'b101001001;
				8'b1010101: c <= 9'b110001100;
				8'b111011: c <= 9'b1100101;
				8'b1001101: c <= 9'b1100011;
				8'b111111: c <= 9'b100000001;
				8'b1101110: c <= 9'b1111001;
				8'b1111011: c <= 9'b100101001;
				8'b1001011: c <= 9'b1110111;
				8'b1101111: c <= 9'b1001100;
				8'b1101000: c <= 9'b110101110;
				8'b101100: c <= 9'b111000101;
				8'b100100: c <= 9'b1010110;
				8'b1111000: c <= 9'b101000111;
				8'b1000101: c <= 9'b111001000;
				8'b1011001: c <= 9'b111111001;
				8'b110100: c <= 9'b1111000;
				8'b1111001: c <= 9'b101010011;
				8'b1110001: c <= 9'b1001010;
				8'b1001111: c <= 9'b100000000;
				8'b1100101: c <= 9'b10001101;
				8'b1111110: c <= 9'b111111110;
				8'b1111100: c <= 9'b110111110;
				8'b1010110: c <= 9'b100010111;
				8'b110010: c <= 9'b11110100;
				8'b1101101: c <= 9'b10101101;
				8'b100011: c <= 9'b100001001;
				8'b1110101: c <= 9'b101010110;
				8'b1111101: c <= 9'b100110;
				8'b101001: c <= 9'b101001001;
				8'b1010010: c <= 9'b111000101;
				8'b1011000: c <= 9'b1100011;
				8'b101110: c <= 9'b11101100;
				8'b1000001: c <= 9'b11101;
				default: c <= 9'b0;
			endcase
			9'b100011010 : case(di)
				8'b1000011: c <= 9'b100001100;
				8'b101000: c <= 9'b100110010;
				8'b111010: c <= 9'b111011011;
				8'b110110: c <= 9'b11001101;
				8'b1100100: c <= 9'b110001100;
				8'b1000000: c <= 9'b101011101;
				8'b1110110: c <= 9'b110101100;
				8'b100101: c <= 9'b10100101;
				8'b101111: c <= 9'b111111011;
				8'b100110: c <= 9'b11001101;
				8'b1100011: c <= 9'b100000000;
				8'b1001000: c <= 9'b110001101;
				8'b111000: c <= 9'b11000111;
				8'b110001: c <= 9'b100110100;
				8'b1010111: c <= 9'b1010001;
				8'b1001110: c <= 9'b110010100;
				8'b1101010: c <= 9'b100111010;
				8'b1001001: c <= 9'b110000101;
				8'b1100000: c <= 9'b100010001;
				8'b110111: c <= 9'b11110101;
				8'b1011101: c <= 9'b110100010;
				8'b1011011: c <= 9'b100011101;
				8'b111001: c <= 9'b1010000;
				8'b1001010: c <= 9'b10011101;
				8'b110011: c <= 9'b11011000;
				8'b1101100: c <= 9'b101011111;
				8'b1110111: c <= 9'b111100111;
				8'b101011: c <= 9'b110000011;
				8'b1101011: c <= 9'b110010010;
				8'b111100: c <= 9'b110000010;
				8'b1000111: c <= 9'b10010000;
				8'b1011111: c <= 9'b1111101;
				8'b1110100: c <= 9'b110101011;
				8'b101101: c <= 9'b110110110;
				8'b1010011: c <= 9'b110001000;
				8'b1100001: c <= 9'b10111101;
				8'b110101: c <= 9'b100111011;
				8'b1000100: c <= 9'b11011110;
				8'b1010001: c <= 9'b100101110;
				8'b1010100: c <= 9'b1000101;
				8'b1100110: c <= 9'b110001000;
				8'b101010: c <= 9'b1110111;
				8'b1011110: c <= 9'b110101010;
				8'b1100111: c <= 9'b11010100;
				8'b1011010: c <= 9'b110011011;
				8'b1000010: c <= 9'b1011000;
				8'b111101: c <= 9'b1111011;
				8'b110000: c <= 9'b101011000;
				8'b111110: c <= 9'b111000111;
				8'b1100010: c <= 9'b111101100;
				8'b1110000: c <= 9'b11010100;
				8'b1101001: c <= 9'b1111111;
				8'b1110011: c <= 9'b10111001;
				8'b1001100: c <= 9'b11010011;
				8'b100001: c <= 9'b101101010;
				8'b1000110: c <= 9'b10000001;
				8'b1110010: c <= 9'b101101;
				8'b1010000: c <= 9'b111111011;
				8'b1111010: c <= 9'b11001000;
				8'b1010101: c <= 9'b1000000;
				8'b111011: c <= 9'b11100001;
				8'b1001101: c <= 9'b1110100;
				8'b111111: c <= 9'b10101110;
				8'b1101110: c <= 9'b111;
				8'b1111011: c <= 9'b100111101;
				8'b1001011: c <= 9'b11101;
				8'b1101111: c <= 9'b110011;
				8'b1101000: c <= 9'b111011011;
				8'b101100: c <= 9'b1010010;
				8'b100100: c <= 9'b100010111;
				8'b1111000: c <= 9'b100011100;
				8'b1000101: c <= 9'b1110000;
				8'b1011001: c <= 9'b110000110;
				8'b110100: c <= 9'b111110101;
				8'b1111001: c <= 9'b110000010;
				8'b1110001: c <= 9'b1100101;
				8'b1001111: c <= 9'b100001100;
				8'b1100101: c <= 9'b110011101;
				8'b1111110: c <= 9'b10001111;
				8'b1111100: c <= 9'b10101100;
				8'b1010110: c <= 9'b1001001;
				8'b110010: c <= 9'b110100100;
				8'b1101101: c <= 9'b1010111;
				8'b100011: c <= 9'b110100010;
				8'b1110101: c <= 9'b1111010;
				8'b1111101: c <= 9'b101101;
				8'b101001: c <= 9'b10010100;
				8'b1010010: c <= 9'b111111000;
				8'b1011000: c <= 9'b10000011;
				8'b101110: c <= 9'b100011101;
				8'b1000001: c <= 9'b1001110;
				default: c <= 9'b0;
			endcase
			9'b10101101 : case(di)
				8'b1000011: c <= 9'b11100001;
				8'b101000: c <= 9'b101101011;
				8'b111010: c <= 9'b10000110;
				8'b110110: c <= 9'b11011001;
				8'b1100100: c <= 9'b100110100;
				8'b1000000: c <= 9'b11110;
				8'b1110110: c <= 9'b10111001;
				8'b100101: c <= 9'b101101;
				8'b101111: c <= 9'b11011110;
				8'b100110: c <= 9'b10111000;
				8'b1100011: c <= 9'b1010111;
				8'b1001000: c <= 9'b11111;
				8'b111000: c <= 9'b110101100;
				8'b110001: c <= 9'b10111011;
				8'b1010111: c <= 9'b11110011;
				8'b1001110: c <= 9'b101011110;
				8'b1101010: c <= 9'b11000100;
				8'b1001001: c <= 9'b11001010;
				8'b1100000: c <= 9'b10001110;
				8'b110111: c <= 9'b10010001;
				8'b1011101: c <= 9'b10101011;
				8'b1011011: c <= 9'b101011011;
				8'b111001: c <= 9'b10000101;
				8'b1001010: c <= 9'b10110;
				8'b110011: c <= 9'b100101010;
				8'b1101100: c <= 9'b101001011;
				8'b1110111: c <= 9'b111010110;
				8'b101011: c <= 9'b110101;
				8'b1101011: c <= 9'b111010110;
				8'b111100: c <= 9'b100010000;
				8'b1000111: c <= 9'b101110010;
				8'b1011111: c <= 9'b10111001;
				8'b1110100: c <= 9'b11001;
				8'b101101: c <= 9'b1101010;
				8'b1010011: c <= 9'b111000;
				8'b1100001: c <= 9'b110001010;
				8'b110101: c <= 9'b100000101;
				8'b1000100: c <= 9'b11110111;
				8'b1010001: c <= 9'b111011011;
				8'b1010100: c <= 9'b100011100;
				8'b1100110: c <= 9'b100111101;
				8'b101010: c <= 9'b101011101;
				8'b1011110: c <= 9'b111000000;
				8'b1100111: c <= 9'b11000100;
				8'b1011010: c <= 9'b101111000;
				8'b1000010: c <= 9'b10110011;
				8'b111101: c <= 9'b110111;
				8'b110000: c <= 9'b100110000;
				8'b111110: c <= 9'b10011000;
				8'b1100010: c <= 9'b1000101;
				8'b1110000: c <= 9'b101001110;
				8'b1101001: c <= 9'b111000100;
				8'b1110011: c <= 9'b11111000;
				8'b1001100: c <= 9'b11100;
				8'b100001: c <= 9'b100000100;
				8'b1000110: c <= 9'b11011110;
				8'b1110010: c <= 9'b110011110;
				8'b1010000: c <= 9'b11001000;
				8'b1111010: c <= 9'b11110111;
				8'b1010101: c <= 9'b10011;
				8'b111011: c <= 9'b1100001;
				8'b1001101: c <= 9'b101000;
				8'b111111: c <= 9'b101101101;
				8'b1101110: c <= 9'b11010101;
				8'b1111011: c <= 9'b1000101;
				8'b1001011: c <= 9'b110110110;
				8'b1101111: c <= 9'b10100111;
				8'b1101000: c <= 9'b10111001;
				8'b101100: c <= 9'b100010110;
				8'b100100: c <= 9'b110011110;
				8'b1111000: c <= 9'b101010000;
				8'b1000101: c <= 9'b110101110;
				8'b1011001: c <= 9'b111000101;
				8'b110100: c <= 9'b101110110;
				8'b1111001: c <= 9'b101100001;
				8'b1110001: c <= 9'b111111101;
				8'b1001111: c <= 9'b1000000;
				8'b1100101: c <= 9'b1100000;
				8'b1111110: c <= 9'b111100111;
				8'b1111100: c <= 9'b10110100;
				8'b1010110: c <= 9'b10001011;
				8'b110010: c <= 9'b110101111;
				8'b1101101: c <= 9'b1001101;
				8'b100011: c <= 9'b1001;
				8'b1110101: c <= 9'b1010011;
				8'b1111101: c <= 9'b1110000;
				8'b101001: c <= 9'b1111110;
				8'b1010010: c <= 9'b110100111;
				8'b1011000: c <= 9'b111010110;
				8'b101110: c <= 9'b110101101;
				8'b1000001: c <= 9'b100011111;
				default: c <= 9'b0;
			endcase
			9'b10000111 : case(di)
				8'b1000011: c <= 9'b111101001;
				8'b101000: c <= 9'b110000;
				8'b111010: c <= 9'b101000011;
				8'b110110: c <= 9'b101101;
				8'b1100100: c <= 9'b101001110;
				8'b1000000: c <= 9'b111011001;
				8'b1110110: c <= 9'b11011110;
				8'b100101: c <= 9'b1111100;
				8'b101111: c <= 9'b11110011;
				8'b100110: c <= 9'b111101101;
				8'b1100011: c <= 9'b10001111;
				8'b1001000: c <= 9'b110000;
				8'b111000: c <= 9'b10010001;
				8'b110001: c <= 9'b11001111;
				8'b1010111: c <= 9'b100011111;
				8'b1001110: c <= 9'b10;
				8'b1101010: c <= 9'b10100000;
				8'b1001001: c <= 9'b100010010;
				8'b1100000: c <= 9'b111000010;
				8'b110111: c <= 9'b11011110;
				8'b1011101: c <= 9'b111110000;
				8'b1011011: c <= 9'b1000001;
				8'b111001: c <= 9'b111101101;
				8'b1001010: c <= 9'b10101101;
				8'b110011: c <= 9'b11111100;
				8'b1101100: c <= 9'b101101;
				8'b1110111: c <= 9'b110001010;
				8'b101011: c <= 9'b10111;
				8'b1101011: c <= 9'b101011101;
				8'b111100: c <= 9'b10011011;
				8'b1000111: c <= 9'b110100;
				8'b1011111: c <= 9'b100100010;
				8'b1110100: c <= 9'b110101;
				8'b101101: c <= 9'b111100;
				8'b1010011: c <= 9'b1011100;
				8'b1100001: c <= 9'b111111110;
				8'b110101: c <= 9'b11111010;
				8'b1000100: c <= 9'b111011011;
				8'b1010001: c <= 9'b111010110;
				8'b1010100: c <= 9'b101101010;
				8'b1100110: c <= 9'b100001011;
				8'b101010: c <= 9'b100010110;
				8'b1011110: c <= 9'b101110010;
				8'b1100111: c <= 9'b110000001;
				8'b1011010: c <= 9'b10111111;
				8'b1000010: c <= 9'b101000111;
				8'b111101: c <= 9'b100111000;
				8'b110000: c <= 9'b111111011;
				8'b111110: c <= 9'b1011011;
				8'b1100010: c <= 9'b10101111;
				8'b1110000: c <= 9'b10110100;
				8'b1101001: c <= 9'b11111000;
				8'b1110011: c <= 9'b10110010;
				8'b1001100: c <= 9'b111100;
				8'b100001: c <= 9'b100001101;
				8'b1000110: c <= 9'b1100101;
				8'b1110010: c <= 9'b100001100;
				8'b1010000: c <= 9'b101110;
				8'b1111010: c <= 9'b11110;
				8'b1010101: c <= 9'b101100;
				8'b111011: c <= 9'b11011110;
				8'b1001101: c <= 9'b100111010;
				8'b111111: c <= 9'b11010100;
				8'b1101110: c <= 9'b100001010;
				8'b1111011: c <= 9'b101111000;
				8'b1001011: c <= 9'b11101111;
				8'b1101111: c <= 9'b100010100;
				8'b1101000: c <= 9'b10101111;
				8'b101100: c <= 9'b100011111;
				8'b100100: c <= 9'b110;
				8'b1111000: c <= 9'b10110011;
				8'b1000101: c <= 9'b11111;
				8'b1011001: c <= 9'b110001001;
				8'b110100: c <= 9'b101000101;
				8'b1111001: c <= 9'b10101001;
				8'b1110001: c <= 9'b110100111;
				8'b1001111: c <= 9'b111000100;
				8'b1100101: c <= 9'b111001110;
				8'b1111110: c <= 9'b100101110;
				8'b1111100: c <= 9'b1001001;
				8'b1010110: c <= 9'b100101010;
				8'b110010: c <= 9'b111111011;
				8'b1101101: c <= 9'b11111;
				8'b100011: c <= 9'b110100100;
				8'b1110101: c <= 9'b101001010;
				8'b1111101: c <= 9'b1100110;
				8'b101001: c <= 9'b10111100;
				8'b1010010: c <= 9'b110010001;
				8'b1011000: c <= 9'b10011;
				8'b101110: c <= 9'b10111100;
				8'b1000001: c <= 9'b101110110;
				default: c <= 9'b0;
			endcase
			9'b101000001 : case(di)
				8'b1000011: c <= 9'b1001010;
				8'b101000: c <= 9'b111111011;
				8'b111010: c <= 9'b1010101;
				8'b110110: c <= 9'b11110010;
				8'b1100100: c <= 9'b100000000;
				8'b1000000: c <= 9'b10001101;
				8'b1110110: c <= 9'b1100100;
				8'b100101: c <= 9'b11100011;
				8'b101111: c <= 9'b1000;
				8'b100110: c <= 9'b101011000;
				8'b1100011: c <= 9'b101001010;
				8'b1001000: c <= 9'b11010000;
				8'b111000: c <= 9'b11000011;
				8'b110001: c <= 9'b100000110;
				8'b1010111: c <= 9'b10011000;
				8'b1001110: c <= 9'b1001101;
				8'b1101010: c <= 9'b101111001;
				8'b1001001: c <= 9'b10010110;
				8'b1100000: c <= 9'b100110100;
				8'b110111: c <= 9'b110111111;
				8'b1011101: c <= 9'b11111110;
				8'b1011011: c <= 9'b100001011;
				8'b111001: c <= 9'b111100000;
				8'b1001010: c <= 9'b111000101;
				8'b110011: c <= 9'b111100;
				8'b1101100: c <= 9'b101100010;
				8'b1110111: c <= 9'b100100111;
				8'b101011: c <= 9'b100111010;
				8'b1101011: c <= 9'b111100111;
				8'b111100: c <= 9'b11110011;
				8'b1000111: c <= 9'b101110011;
				8'b1011111: c <= 9'b101011010;
				8'b1110100: c <= 9'b10011;
				8'b101101: c <= 9'b111111000;
				8'b1010011: c <= 9'b10001110;
				8'b1100001: c <= 9'b100101;
				8'b110101: c <= 9'b111011010;
				8'b1000100: c <= 9'b10101010;
				8'b1010001: c <= 9'b11111000;
				8'b1010100: c <= 9'b10110001;
				8'b1100110: c <= 9'b101010011;
				8'b101010: c <= 9'b100110101;
				8'b1011110: c <= 9'b101;
				8'b1100111: c <= 9'b110001;
				8'b1011010: c <= 9'b10010011;
				8'b1000010: c <= 9'b101010011;
				8'b111101: c <= 9'b101001111;
				8'b110000: c <= 9'b100111001;
				8'b111110: c <= 9'b11100001;
				8'b1100010: c <= 9'b1000110;
				8'b1110000: c <= 9'b11111100;
				8'b1101001: c <= 9'b10101100;
				8'b1110011: c <= 9'b111001101;
				8'b1001100: c <= 9'b100111010;
				8'b100001: c <= 9'b100010010;
				8'b1000110: c <= 9'b101000;
				8'b1110010: c <= 9'b101011101;
				8'b1010000: c <= 9'b110110110;
				8'b1111010: c <= 9'b11011100;
				8'b1010101: c <= 9'b110001011;
				8'b111011: c <= 9'b11111101;
				8'b1001101: c <= 9'b100101010;
				8'b111111: c <= 9'b11001011;
				8'b1101110: c <= 9'b11000111;
				8'b1111011: c <= 9'b100000110;
				8'b1001011: c <= 9'b101001011;
				8'b1101111: c <= 9'b111111101;
				8'b1101000: c <= 9'b110101001;
				8'b101100: c <= 9'b101100100;
				8'b100100: c <= 9'b100100111;
				8'b1111000: c <= 9'b111111011;
				8'b1000101: c <= 9'b10000111;
				8'b1011001: c <= 9'b11000110;
				8'b110100: c <= 9'b111100010;
				8'b1111001: c <= 9'b10010011;
				8'b1110001: c <= 9'b101010101;
				8'b1001111: c <= 9'b100010111;
				8'b1100101: c <= 9'b11111110;
				8'b1111110: c <= 9'b10010100;
				8'b1111100: c <= 9'b100011000;
				8'b1010110: c <= 9'b101111000;
				8'b110010: c <= 9'b100101010;
				8'b1101101: c <= 9'b111000101;
				8'b100011: c <= 9'b111;
				8'b1110101: c <= 9'b100110110;
				8'b1111101: c <= 9'b100000000;
				8'b101001: c <= 9'b10111110;
				8'b1010010: c <= 9'b111101;
				8'b1011000: c <= 9'b10000000;
				8'b101110: c <= 9'b100100010;
				8'b1000001: c <= 9'b101100110;
				default: c <= 9'b0;
			endcase
			9'b101011111 : case(di)
				8'b1000011: c <= 9'b100010;
				8'b101000: c <= 9'b10110111;
				8'b111010: c <= 9'b11110010;
				8'b110110: c <= 9'b11000010;
				8'b1100100: c <= 9'b101001010;
				8'b1000000: c <= 9'b101011;
				8'b1110110: c <= 9'b101010010;
				8'b100101: c <= 9'b10101010;
				8'b101111: c <= 9'b1011;
				8'b100110: c <= 9'b111101000;
				8'b1100011: c <= 9'b11011010;
				8'b1001000: c <= 9'b111101;
				8'b111000: c <= 9'b10010110;
				8'b110001: c <= 9'b1100111;
				8'b1010111: c <= 9'b100001010;
				8'b1001110: c <= 9'b111111001;
				8'b1101010: c <= 9'b11011;
				8'b1001001: c <= 9'b100001;
				8'b1100000: c <= 9'b100010101;
				8'b110111: c <= 9'b10100;
				8'b1011101: c <= 9'b11101101;
				8'b1011011: c <= 9'b111001000;
				8'b111001: c <= 9'b110011101;
				8'b1001010: c <= 9'b111010100;
				8'b110011: c <= 9'b110010011;
				8'b1101100: c <= 9'b101011011;
				8'b1110111: c <= 9'b100111;
				8'b101011: c <= 9'b100100101;
				8'b1101011: c <= 9'b100100111;
				8'b111100: c <= 9'b11001110;
				8'b1000111: c <= 9'b100111001;
				8'b1011111: c <= 9'b10100100;
				8'b1110100: c <= 9'b111000011;
				8'b101101: c <= 9'b110001100;
				8'b1010011: c <= 9'b111100000;
				8'b1100001: c <= 9'b100110011;
				8'b110101: c <= 9'b11001000;
				8'b1000100: c <= 9'b1000011;
				8'b1010001: c <= 9'b11011010;
				8'b1010100: c <= 9'b101010110;
				8'b1100110: c <= 9'b111110001;
				8'b101010: c <= 9'b110011011;
				8'b1011110: c <= 9'b111001;
				8'b1100111: c <= 9'b110110000;
				8'b1011010: c <= 9'b101110001;
				8'b1000010: c <= 9'b110110101;
				8'b111101: c <= 9'b110101011;
				8'b110000: c <= 9'b111001011;
				8'b111110: c <= 9'b10101001;
				8'b1100010: c <= 9'b100101000;
				8'b1110000: c <= 9'b1000;
				8'b1101001: c <= 9'b101000110;
				8'b1110011: c <= 9'b101100111;
				8'b1001100: c <= 9'b111100100;
				8'b100001: c <= 9'b111101111;
				8'b1000110: c <= 9'b111001010;
				8'b1110010: c <= 9'b10011111;
				8'b1010000: c <= 9'b110011000;
				8'b1111010: c <= 9'b1010101;
				8'b1010101: c <= 9'b11111101;
				8'b111011: c <= 9'b1011011;
				8'b1001101: c <= 9'b111111110;
				8'b111111: c <= 9'b1100010;
				8'b1101110: c <= 9'b11110110;
				8'b1111011: c <= 9'b100101010;
				8'b1001011: c <= 9'b110010111;
				8'b1101111: c <= 9'b101110011;
				8'b1101000: c <= 9'b100101001;
				8'b101100: c <= 9'b10100000;
				8'b100100: c <= 9'b100111101;
				8'b1111000: c <= 9'b100110000;
				8'b1000101: c <= 9'b110000000;
				8'b1011001: c <= 9'b11010101;
				8'b110100: c <= 9'b111010111;
				8'b1111001: c <= 9'b110010101;
				8'b1110001: c <= 9'b101100001;
				8'b1001111: c <= 9'b101010;
				8'b1100101: c <= 9'b101101111;
				8'b1111110: c <= 9'b10010001;
				8'b1111100: c <= 9'b101001100;
				8'b1010110: c <= 9'b1001010;
				8'b110010: c <= 9'b11100111;
				8'b1101101: c <= 9'b110101010;
				8'b100011: c <= 9'b10111010;
				8'b1110101: c <= 9'b10100011;
				8'b1111101: c <= 9'b111;
				8'b101001: c <= 9'b1001011;
				8'b1010010: c <= 9'b100100111;
				8'b1011000: c <= 9'b1100100;
				8'b101110: c <= 9'b111111101;
				8'b1000001: c <= 9'b1011110;
				default: c <= 9'b0;
			endcase
			9'b10000001 : case(di)
				8'b1000011: c <= 9'b11001100;
				8'b101000: c <= 9'b101011011;
				8'b111010: c <= 9'b101010010;
				8'b110110: c <= 9'b110101001;
				8'b1100100: c <= 9'b1100111;
				8'b1000000: c <= 9'b10101011;
				8'b1110110: c <= 9'b11010100;
				8'b100101: c <= 9'b11110001;
				8'b101111: c <= 9'b111100110;
				8'b100110: c <= 9'b110010101;
				8'b1100011: c <= 9'b101000110;
				8'b1001000: c <= 9'b11001100;
				8'b111000: c <= 9'b111001100;
				8'b110001: c <= 9'b111100011;
				8'b1010111: c <= 9'b110011110;
				8'b1001110: c <= 9'b11011110;
				8'b1101010: c <= 9'b101000010;
				8'b1001001: c <= 9'b10110;
				8'b1100000: c <= 9'b101001110;
				8'b110111: c <= 9'b11001000;
				8'b1011101: c <= 9'b1111100;
				8'b1011011: c <= 9'b10001110;
				8'b111001: c <= 9'b10110100;
				8'b1001010: c <= 9'b11010100;
				8'b110011: c <= 9'b11;
				8'b1101100: c <= 9'b101111001;
				8'b1110111: c <= 9'b10001001;
				8'b101011: c <= 9'b110110011;
				8'b1101011: c <= 9'b10101110;
				8'b111100: c <= 9'b1111100;
				8'b1000111: c <= 9'b11001100;
				8'b1011111: c <= 9'b111110101;
				8'b1110100: c <= 9'b100110100;
				8'b101101: c <= 9'b110101100;
				8'b1010011: c <= 9'b100001110;
				8'b1100001: c <= 9'b10001100;
				8'b110101: c <= 9'b101101101;
				8'b1000100: c <= 9'b11100010;
				8'b1010001: c <= 9'b11000010;
				8'b1010100: c <= 9'b100011001;
				8'b1100110: c <= 9'b100001110;
				8'b101010: c <= 9'b111001011;
				8'b1011110: c <= 9'b110110011;
				8'b1100111: c <= 9'b110100;
				8'b1011010: c <= 9'b101010101;
				8'b1000010: c <= 9'b10001011;
				8'b111101: c <= 9'b111001011;
				8'b110000: c <= 9'b10001100;
				8'b111110: c <= 9'b110100001;
				8'b1100010: c <= 9'b111100001;
				8'b1110000: c <= 9'b100111111;
				8'b1101001: c <= 9'b100111010;
				8'b1110011: c <= 9'b110000;
				8'b1001100: c <= 9'b110111;
				8'b100001: c <= 9'b111001010;
				8'b1000110: c <= 9'b111000011;
				8'b1110010: c <= 9'b101111110;
				8'b1010000: c <= 9'b110001011;
				8'b1111010: c <= 9'b1000111;
				8'b1010101: c <= 9'b111100100;
				8'b111011: c <= 9'b111010111;
				8'b1001101: c <= 9'b101110111;
				8'b111111: c <= 9'b100010101;
				8'b1101110: c <= 9'b110111111;
				8'b1111011: c <= 9'b110110010;
				8'b1001011: c <= 9'b111001100;
				8'b1101111: c <= 9'b101001001;
				8'b1101000: c <= 9'b101010011;
				8'b101100: c <= 9'b111111101;
				8'b100100: c <= 9'b101101110;
				8'b1111000: c <= 9'b10111;
				8'b1000101: c <= 9'b110101;
				8'b1011001: c <= 9'b110100100;
				8'b110100: c <= 9'b100111011;
				8'b1111001: c <= 9'b100011101;
				8'b1110001: c <= 9'b100010111;
				8'b1001111: c <= 9'b101010101;
				8'b1100101: c <= 9'b101101011;
				8'b1111110: c <= 9'b1100100;
				8'b1111100: c <= 9'b100111000;
				8'b1010110: c <= 9'b10010011;
				8'b110010: c <= 9'b11011110;
				8'b1101101: c <= 9'b110100111;
				8'b100011: c <= 9'b1001011;
				8'b1110101: c <= 9'b111111000;
				8'b1111101: c <= 9'b111111000;
				8'b101001: c <= 9'b100111100;
				8'b1010010: c <= 9'b111100;
				8'b1011000: c <= 9'b111100;
				8'b101110: c <= 9'b10011001;
				8'b1000001: c <= 9'b1011110;
				default: c <= 9'b0;
			endcase
			9'b110110111 : case(di)
				8'b1000011: c <= 9'b110101011;
				8'b101000: c <= 9'b111001110;
				8'b111010: c <= 9'b111000;
				8'b110110: c <= 9'b11000001;
				8'b1100100: c <= 9'b10011;
				8'b1000000: c <= 9'b1111100;
				8'b1110110: c <= 9'b101100011;
				8'b100101: c <= 9'b1100000;
				8'b101111: c <= 9'b1001001;
				8'b100110: c <= 9'b100111011;
				8'b1100011: c <= 9'b101100101;
				8'b1001000: c <= 9'b110010010;
				8'b111000: c <= 9'b101011000;
				8'b110001: c <= 9'b111010110;
				8'b1010111: c <= 9'b110110011;
				8'b1001110: c <= 9'b100010110;
				8'b1101010: c <= 9'b111010111;
				8'b1001001: c <= 9'b1101110;
				8'b1100000: c <= 9'b11110110;
				8'b110111: c <= 9'b110100111;
				8'b1011101: c <= 9'b101001001;
				8'b1011011: c <= 9'b11000111;
				8'b111001: c <= 9'b100;
				8'b1001010: c <= 9'b110110;
				8'b110011: c <= 9'b101001;
				8'b1101100: c <= 9'b111001010;
				8'b1110111: c <= 9'b100001001;
				8'b101011: c <= 9'b100101000;
				8'b1101011: c <= 9'b101100001;
				8'b111100: c <= 9'b11101001;
				8'b1000111: c <= 9'b111100010;
				8'b1011111: c <= 9'b100110011;
				8'b1110100: c <= 9'b110011;
				8'b101101: c <= 9'b101010;
				8'b1010011: c <= 9'b100001110;
				8'b1100001: c <= 9'b10011011;
				8'b110101: c <= 9'b11100110;
				8'b1000100: c <= 9'b10100;
				8'b1010001: c <= 9'b10000010;
				8'b1010100: c <= 9'b100111011;
				8'b1100110: c <= 9'b111101001;
				8'b101010: c <= 9'b110011011;
				8'b1011110: c <= 9'b10000111;
				8'b1100111: c <= 9'b101010001;
				8'b1011010: c <= 9'b111010000;
				8'b1000010: c <= 9'b110000110;
				8'b111101: c <= 9'b1101001;
				8'b110000: c <= 9'b111000100;
				8'b111110: c <= 9'b1001110;
				8'b1100010: c <= 9'b100110011;
				8'b1110000: c <= 9'b100111000;
				8'b1101001: c <= 9'b1110000;
				8'b1110011: c <= 9'b101111001;
				8'b1001100: c <= 9'b100101010;
				8'b100001: c <= 9'b10011001;
				8'b1000110: c <= 9'b100010100;
				8'b1110010: c <= 9'b11100011;
				8'b1010000: c <= 9'b111011101;
				8'b1111010: c <= 9'b111101;
				8'b1010101: c <= 9'b1110100;
				8'b111011: c <= 9'b111010100;
				8'b1001101: c <= 9'b10010000;
				8'b111111: c <= 9'b100001001;
				8'b1101110: c <= 9'b10101001;
				8'b1111011: c <= 9'b11111;
				8'b1001011: c <= 9'b11001110;
				8'b1101111: c <= 9'b100100110;
				8'b1101000: c <= 9'b1000011;
				8'b101100: c <= 9'b111011;
				8'b100100: c <= 9'b1011110;
				8'b1111000: c <= 9'b110110110;
				8'b1000101: c <= 9'b10110110;
				8'b1011001: c <= 9'b111101100;
				8'b110100: c <= 9'b1000110;
				8'b1111001: c <= 9'b10110;
				8'b1110001: c <= 9'b111001010;
				8'b1001111: c <= 9'b1111010;
				8'b1100101: c <= 9'b10000;
				8'b1111110: c <= 9'b110011001;
				8'b1111100: c <= 9'b100000111;
				8'b1010110: c <= 9'b1101111;
				8'b110010: c <= 9'b101011000;
				8'b1101101: c <= 9'b101000001;
				8'b100011: c <= 9'b111101010;
				8'b1110101: c <= 9'b1100111;
				8'b1111101: c <= 9'b111101110;
				8'b101001: c <= 9'b1101001;
				8'b1010010: c <= 9'b110010111;
				8'b1011000: c <= 9'b1010010;
				8'b101110: c <= 9'b1111001;
				8'b1000001: c <= 9'b110001001;
				default: c <= 9'b0;
			endcase
			9'b100101011 : case(di)
				8'b1000011: c <= 9'b10100100;
				8'b101000: c <= 9'b10111110;
				8'b111010: c <= 9'b110001101;
				8'b110110: c <= 9'b101111111;
				8'b1100100: c <= 9'b100101111;
				8'b1000000: c <= 9'b10100011;
				8'b1110110: c <= 9'b10101011;
				8'b100101: c <= 9'b111100100;
				8'b101111: c <= 9'b1100000;
				8'b100110: c <= 9'b110010100;
				8'b1100011: c <= 9'b11010001;
				8'b1001000: c <= 9'b1001;
				8'b111000: c <= 9'b111001100;
				8'b110001: c <= 9'b11011001;
				8'b1010111: c <= 9'b101000;
				8'b1001110: c <= 9'b110110100;
				8'b1101010: c <= 9'b110;
				8'b1001001: c <= 9'b111111000;
				8'b1100000: c <= 9'b101100110;
				8'b110111: c <= 9'b110011010;
				8'b1011101: c <= 9'b100110010;
				8'b1011011: c <= 9'b1;
				8'b111001: c <= 9'b110111001;
				8'b1001010: c <= 9'b1111011;
				8'b110011: c <= 9'b110101;
				8'b1101100: c <= 9'b1001011;
				8'b1110111: c <= 9'b11110001;
				8'b101011: c <= 9'b11001011;
				8'b1101011: c <= 9'b100101111;
				8'b111100: c <= 9'b110101010;
				8'b1000111: c <= 9'b100001;
				8'b1011111: c <= 9'b101011110;
				8'b1110100: c <= 9'b111100011;
				8'b101101: c <= 9'b10000000;
				8'b1010011: c <= 9'b110110011;
				8'b1100001: c <= 9'b1011100;
				8'b110101: c <= 9'b11010010;
				8'b1000100: c <= 9'b11110001;
				8'b1010001: c <= 9'b10011001;
				8'b1010100: c <= 9'b101010110;
				8'b1100110: c <= 9'b100111110;
				8'b101010: c <= 9'b10100111;
				8'b1011110: c <= 9'b110101100;
				8'b1100111: c <= 9'b110001;
				8'b1011010: c <= 9'b11001000;
				8'b1000010: c <= 9'b110001010;
				8'b111101: c <= 9'b1000010;
				8'b110000: c <= 9'b111001100;
				8'b111110: c <= 9'b1001100;
				8'b1100010: c <= 9'b11110111;
				8'b1110000: c <= 9'b100010001;
				8'b1101001: c <= 9'b10100010;
				8'b1110011: c <= 9'b1010010;
				8'b1001100: c <= 9'b11111001;
				8'b100001: c <= 9'b1100110;
				8'b1000110: c <= 9'b10;
				8'b1110010: c <= 9'b111101110;
				8'b1010000: c <= 9'b1110101;
				8'b1111010: c <= 9'b110111011;
				8'b1010101: c <= 9'b111010000;
				8'b111011: c <= 9'b111010;
				8'b1001101: c <= 9'b101111000;
				8'b111111: c <= 9'b101110;
				8'b1101110: c <= 9'b111110011;
				8'b1111011: c <= 9'b1001010;
				8'b1001011: c <= 9'b101110100;
				8'b1101111: c <= 9'b11000;
				8'b1101000: c <= 9'b110011010;
				8'b101100: c <= 9'b11110100;
				8'b100100: c <= 9'b10;
				8'b1111000: c <= 9'b101011110;
				8'b1000101: c <= 9'b110111010;
				8'b1011001: c <= 9'b111100011;
				8'b110100: c <= 9'b110100000;
				8'b1111001: c <= 9'b1010011;
				8'b1110001: c <= 9'b111001000;
				8'b1001111: c <= 9'b111111101;
				8'b1100101: c <= 9'b10111001;
				8'b1111110: c <= 9'b11111000;
				8'b1111100: c <= 9'b100010101;
				8'b1010110: c <= 9'b110010101;
				8'b110010: c <= 9'b101101100;
				8'b1101101: c <= 9'b111101;
				8'b100011: c <= 9'b101110000;
				8'b1110101: c <= 9'b100111010;
				8'b1111101: c <= 9'b110010;
				8'b101001: c <= 9'b111100001;
				8'b1010010: c <= 9'b1111011;
				8'b1011000: c <= 9'b11011010;
				8'b101110: c <= 9'b11101011;
				8'b1000001: c <= 9'b101100100;
				default: c <= 9'b0;
			endcase
			9'b110010001 : case(di)
				8'b1000011: c <= 9'b100011000;
				8'b101000: c <= 9'b11110010;
				8'b111010: c <= 9'b100111111;
				8'b110110: c <= 9'b10010110;
				8'b1100100: c <= 9'b110101011;
				8'b1000000: c <= 9'b11111001;
				8'b1110110: c <= 9'b11110100;
				8'b100101: c <= 9'b110111000;
				8'b101111: c <= 9'b10111011;
				8'b100110: c <= 9'b101010;
				8'b1100011: c <= 9'b100111111;
				8'b1001000: c <= 9'b10101010;
				8'b111000: c <= 9'b110101101;
				8'b110001: c <= 9'b100110110;
				8'b1010111: c <= 9'b1010000;
				8'b1001110: c <= 9'b11000001;
				8'b1101010: c <= 9'b101000011;
				8'b1001001: c <= 9'b101101010;
				8'b1100000: c <= 9'b110100;
				8'b110111: c <= 9'b110111001;
				8'b1011101: c <= 9'b1011000;
				8'b1011011: c <= 9'b10010100;
				8'b111001: c <= 9'b11101100;
				8'b1001010: c <= 9'b11100;
				8'b110011: c <= 9'b1101101;
				8'b1101100: c <= 9'b110110110;
				8'b1110111: c <= 9'b110000110;
				8'b101011: c <= 9'b11101001;
				8'b1101011: c <= 9'b100100111;
				8'b111100: c <= 9'b100001100;
				8'b1000111: c <= 9'b101100001;
				8'b1011111: c <= 9'b10100111;
				8'b1110100: c <= 9'b111111110;
				8'b101101: c <= 9'b110111110;
				8'b1010011: c <= 9'b100101101;
				8'b1100001: c <= 9'b10001101;
				8'b110101: c <= 9'b1101;
				8'b1000100: c <= 9'b10111110;
				8'b1010001: c <= 9'b100011010;
				8'b1010100: c <= 9'b11000110;
				8'b1100110: c <= 9'b110011011;
				8'b101010: c <= 9'b10100000;
				8'b1011110: c <= 9'b110000;
				8'b1100111: c <= 9'b10100011;
				8'b1011010: c <= 9'b11111;
				8'b1000010: c <= 9'b100100001;
				8'b111101: c <= 9'b100100011;
				8'b110000: c <= 9'b110010;
				8'b111110: c <= 9'b100101101;
				8'b1100010: c <= 9'b1000101;
				8'b1110000: c <= 9'b10101101;
				8'b1101001: c <= 9'b1001100;
				8'b1110011: c <= 9'b10011011;
				8'b1001100: c <= 9'b111000000;
				8'b100001: c <= 9'b111101110;
				8'b1000110: c <= 9'b1000;
				8'b1110010: c <= 9'b110110000;
				8'b1010000: c <= 9'b111110000;
				8'b1111010: c <= 9'b10000110;
				8'b1010101: c <= 9'b100100101;
				8'b111011: c <= 9'b1000010;
				8'b1001101: c <= 9'b100101110;
				8'b111111: c <= 9'b110100101;
				8'b1101110: c <= 9'b111011;
				8'b1111011: c <= 9'b11100110;
				8'b1001011: c <= 9'b110111100;
				8'b1101111: c <= 9'b100011010;
				8'b1101000: c <= 9'b1011011;
				8'b101100: c <= 9'b110101;
				8'b100100: c <= 9'b101001;
				8'b1111000: c <= 9'b100101100;
				8'b1000101: c <= 9'b100010111;
				8'b1011001: c <= 9'b110001101;
				8'b110100: c <= 9'b10100011;
				8'b1111001: c <= 9'b101011000;
				8'b1110001: c <= 9'b1001010;
				8'b1001111: c <= 9'b111000011;
				8'b1100101: c <= 9'b10001101;
				8'b1111110: c <= 9'b11010000;
				8'b1111100: c <= 9'b111101101;
				8'b1010110: c <= 9'b10100100;
				8'b110010: c <= 9'b101010101;
				8'b1101101: c <= 9'b10101110;
				8'b100011: c <= 9'b101100100;
				8'b1110101: c <= 9'b110000001;
				8'b1111101: c <= 9'b11100000;
				8'b101001: c <= 9'b11010011;
				8'b1010010: c <= 9'b10001111;
				8'b1011000: c <= 9'b110001110;
				8'b101110: c <= 9'b110000110;
				8'b1000001: c <= 9'b100001001;
				default: c <= 9'b0;
			endcase
			9'b10001000 : case(di)
				8'b1000011: c <= 9'b1010111;
				8'b101000: c <= 9'b10101100;
				8'b111010: c <= 9'b111010;
				8'b110110: c <= 9'b101000001;
				8'b1100100: c <= 9'b101010011;
				8'b1000000: c <= 9'b100011;
				8'b1110110: c <= 9'b110101110;
				8'b100101: c <= 9'b100010010;
				8'b101111: c <= 9'b11111110;
				8'b100110: c <= 9'b110110011;
				8'b1100011: c <= 9'b101101110;
				8'b1001000: c <= 9'b11010101;
				8'b111000: c <= 9'b110010;
				8'b110001: c <= 9'b1101111;
				8'b1010111: c <= 9'b100010;
				8'b1001110: c <= 9'b1101;
				8'b1101010: c <= 9'b11010000;
				8'b1001001: c <= 9'b10001110;
				8'b1100000: c <= 9'b111010010;
				8'b110111: c <= 9'b100000110;
				8'b1011101: c <= 9'b110000111;
				8'b1011011: c <= 9'b100101110;
				8'b111001: c <= 9'b101011001;
				8'b1001010: c <= 9'b11100010;
				8'b110011: c <= 9'b100111000;
				8'b1101100: c <= 9'b11010;
				8'b1110111: c <= 9'b111110110;
				8'b101011: c <= 9'b10011111;
				8'b1101011: c <= 9'b111110000;
				8'b111100: c <= 9'b100110;
				8'b1000111: c <= 9'b110111010;
				8'b1011111: c <= 9'b111110001;
				8'b1110100: c <= 9'b10011100;
				8'b101101: c <= 9'b101100100;
				8'b1010011: c <= 9'b11001100;
				8'b1100001: c <= 9'b110001000;
				8'b110101: c <= 9'b111110001;
				8'b1000100: c <= 9'b111101000;
				8'b1010001: c <= 9'b11001101;
				8'b1010100: c <= 9'b111111111;
				8'b1100110: c <= 9'b11110010;
				8'b101010: c <= 9'b111011101;
				8'b1011110: c <= 9'b10111010;
				8'b1100111: c <= 9'b110010111;
				8'b1011010: c <= 9'b10110001;
				8'b1000010: c <= 9'b11011100;
				8'b111101: c <= 9'b1100011;
				8'b110000: c <= 9'b111001001;
				8'b111110: c <= 9'b1111101;
				8'b1100010: c <= 9'b100110111;
				8'b1110000: c <= 9'b111100001;
				8'b1101001: c <= 9'b10110001;
				8'b1110011: c <= 9'b10010110;
				8'b1001100: c <= 9'b110111111;
				8'b100001: c <= 9'b1111111;
				8'b1000110: c <= 9'b101100110;
				8'b1110010: c <= 9'b101001111;
				8'b1010000: c <= 9'b110110011;
				8'b1111010: c <= 9'b1101111;
				8'b1010101: c <= 9'b110101101;
				8'b111011: c <= 9'b100000101;
				8'b1001101: c <= 9'b100101110;
				8'b111111: c <= 9'b1111011;
				8'b1101110: c <= 9'b1000001;
				8'b1111011: c <= 9'b10011011;
				8'b1001011: c <= 9'b111111010;
				8'b1101111: c <= 9'b10110010;
				8'b1101000: c <= 9'b11110000;
				8'b101100: c <= 9'b11000010;
				8'b100100: c <= 9'b1101010;
				8'b1111000: c <= 9'b111000000;
				8'b1000101: c <= 9'b10001001;
				8'b1011001: c <= 9'b110111010;
				8'b110100: c <= 9'b110001111;
				8'b1111001: c <= 9'b1000111;
				8'b1110001: c <= 9'b110010010;
				8'b1001111: c <= 9'b100101110;
				8'b1100101: c <= 9'b1110100;
				8'b1111110: c <= 9'b110000010;
				8'b1111100: c <= 9'b101100001;
				8'b1010110: c <= 9'b101111001;
				8'b110010: c <= 9'b101100000;
				8'b1101101: c <= 9'b100011001;
				8'b100011: c <= 9'b1010110;
				8'b1110101: c <= 9'b111100001;
				8'b1111101: c <= 9'b1111100;
				8'b101001: c <= 9'b110111100;
				8'b1010010: c <= 9'b1110010;
				8'b1011000: c <= 9'b100011011;
				8'b101110: c <= 9'b101111010;
				8'b1000001: c <= 9'b101110111;
				default: c <= 9'b0;
			endcase
			9'b100111011 : case(di)
				8'b1000011: c <= 9'b11001010;
				8'b101000: c <= 9'b10101011;
				8'b111010: c <= 9'b10110100;
				8'b110110: c <= 9'b11000010;
				8'b1100100: c <= 9'b1010000;
				8'b1000000: c <= 9'b1001010;
				8'b1110110: c <= 9'b100001100;
				8'b100101: c <= 9'b10001111;
				8'b101111: c <= 9'b100100;
				8'b100110: c <= 9'b101000111;
				8'b1100011: c <= 9'b101011110;
				8'b1001000: c <= 9'b111101010;
				8'b111000: c <= 9'b101100;
				8'b110001: c <= 9'b100111000;
				8'b1010111: c <= 9'b1100110;
				8'b1001110: c <= 9'b11001101;
				8'b1101010: c <= 9'b1000010;
				8'b1001001: c <= 9'b11001111;
				8'b1100000: c <= 9'b11011000;
				8'b110111: c <= 9'b1110111;
				8'b1011101: c <= 9'b100011100;
				8'b1011011: c <= 9'b1010010;
				8'b111001: c <= 9'b100000011;
				8'b1001010: c <= 9'b110101101;
				8'b110011: c <= 9'b100010010;
				8'b1101100: c <= 9'b111100101;
				8'b1110111: c <= 9'b111011011;
				8'b101011: c <= 9'b111111010;
				8'b1101011: c <= 9'b100011001;
				8'b111100: c <= 9'b101000001;
				8'b1000111: c <= 9'b10010011;
				8'b1011111: c <= 9'b100111101;
				8'b1110100: c <= 9'b111100011;
				8'b101101: c <= 9'b100010100;
				8'b1010011: c <= 9'b1011000;
				8'b1100001: c <= 9'b1010111;
				8'b110101: c <= 9'b10;
				8'b1000100: c <= 9'b10000000;
				8'b1010001: c <= 9'b111101000;
				8'b1010100: c <= 9'b10101111;
				8'b1100110: c <= 9'b101110101;
				8'b101010: c <= 9'b110010011;
				8'b1011110: c <= 9'b100001101;
				8'b1100111: c <= 9'b110101;
				8'b1011010: c <= 9'b11100101;
				8'b1000010: c <= 9'b10110110;
				8'b111101: c <= 9'b110010100;
				8'b110000: c <= 9'b100101101;
				8'b111110: c <= 9'b111010111;
				8'b1100010: c <= 9'b10001111;
				8'b1110000: c <= 9'b1110001;
				8'b1101001: c <= 9'b1011100;
				8'b1110011: c <= 9'b1111;
				8'b1001100: c <= 9'b1010111;
				8'b100001: c <= 9'b1000;
				8'b1000110: c <= 9'b101101000;
				8'b1110010: c <= 9'b110111010;
				8'b1010000: c <= 9'b111111011;
				8'b1111010: c <= 9'b10000110;
				8'b1010101: c <= 9'b100100101;
				8'b111011: c <= 9'b110110000;
				8'b1001101: c <= 9'b10011000;
				8'b111111: c <= 9'b10011;
				8'b1101110: c <= 9'b100101010;
				8'b1111011: c <= 9'b10010001;
				8'b1001011: c <= 9'b1001000;
				8'b1101111: c <= 9'b111;
				8'b1101000: c <= 9'b10101;
				8'b101100: c <= 9'b10000011;
				8'b100100: c <= 9'b10000001;
				8'b1111000: c <= 9'b111100001;
				8'b1000101: c <= 9'b1101000;
				8'b1011001: c <= 9'b101100011;
				8'b110100: c <= 9'b101100010;
				8'b1111001: c <= 9'b10100000;
				8'b1110001: c <= 9'b1010010;
				8'b1001111: c <= 9'b1011;
				8'b1100101: c <= 9'b110011100;
				8'b1111110: c <= 9'b110101001;
				8'b1111100: c <= 9'b10011000;
				8'b1010110: c <= 9'b10011100;
				8'b110010: c <= 9'b101101111;
				8'b1101101: c <= 9'b100101110;
				8'b100011: c <= 9'b101001110;
				8'b1110101: c <= 9'b10011111;
				8'b1111101: c <= 9'b1011011;
				8'b101001: c <= 9'b101111010;
				8'b1010010: c <= 9'b101110110;
				8'b1011000: c <= 9'b101110010;
				8'b101110: c <= 9'b1010010;
				8'b1000001: c <= 9'b10001111;
				default: c <= 9'b0;
			endcase
			9'b111010111 : case(di)
				8'b1000011: c <= 9'b101101100;
				8'b101000: c <= 9'b111100001;
				8'b111010: c <= 9'b11100101;
				8'b110110: c <= 9'b1000000;
				8'b1100100: c <= 9'b110100100;
				8'b1000000: c <= 9'b100101110;
				8'b1110110: c <= 9'b111110110;
				8'b100101: c <= 9'b101001010;
				8'b101111: c <= 9'b101011000;
				8'b100110: c <= 9'b110011011;
				8'b1100011: c <= 9'b101010000;
				8'b1001000: c <= 9'b100010001;
				8'b111000: c <= 9'b111000110;
				8'b110001: c <= 9'b10011011;
				8'b1010111: c <= 9'b11100111;
				8'b1001110: c <= 9'b101001110;
				8'b1101010: c <= 9'b101000001;
				8'b1001001: c <= 9'b1011000;
				8'b1100000: c <= 9'b111111011;
				8'b110111: c <= 9'b100011000;
				8'b1011101: c <= 9'b110011111;
				8'b1011011: c <= 9'b110011011;
				8'b111001: c <= 9'b10101;
				8'b1001010: c <= 9'b100101100;
				8'b110011: c <= 9'b1000100;
				8'b1101100: c <= 9'b1001;
				8'b1110111: c <= 9'b10110101;
				8'b101011: c <= 9'b1001100;
				8'b1101011: c <= 9'b10011101;
				8'b111100: c <= 9'b100110;
				8'b1000111: c <= 9'b110110110;
				8'b1011111: c <= 9'b111000101;
				8'b1110100: c <= 9'b101001111;
				8'b101101: c <= 9'b11111110;
				8'b1010011: c <= 9'b11100001;
				8'b1100001: c <= 9'b11010011;
				8'b110101: c <= 9'b100100101;
				8'b1000100: c <= 9'b1011001;
				8'b1010001: c <= 9'b110000;
				8'b1010100: c <= 9'b1101000;
				8'b1100110: c <= 9'b1111;
				8'b101010: c <= 9'b10101001;
				8'b1011110: c <= 9'b101000101;
				8'b1100111: c <= 9'b11100101;
				8'b1011010: c <= 9'b11001101;
				8'b1000010: c <= 9'b101011001;
				8'b111101: c <= 9'b110011100;
				8'b110000: c <= 9'b101101001;
				8'b111110: c <= 9'b101011011;
				8'b1100010: c <= 9'b111001101;
				8'b1110000: c <= 9'b111110001;
				8'b1101001: c <= 9'b100101011;
				8'b1110011: c <= 9'b110010011;
				8'b1001100: c <= 9'b1111100;
				8'b100001: c <= 9'b1001000;
				8'b1000110: c <= 9'b101010010;
				8'b1110010: c <= 9'b10010101;
				8'b1010000: c <= 9'b1101010;
				8'b1111010: c <= 9'b110100111;
				8'b1010101: c <= 9'b100101011;
				8'b111011: c <= 9'b111011;
				8'b1001101: c <= 9'b101000100;
				8'b111111: c <= 9'b11010;
				8'b1101110: c <= 9'b11111100;
				8'b1111011: c <= 9'b101011010;
				8'b1001011: c <= 9'b11001111;
				8'b1101111: c <= 9'b101;
				8'b1101000: c <= 9'b101101011;
				8'b101100: c <= 9'b1001;
				8'b100100: c <= 9'b1000;
				8'b1111000: c <= 9'b100011111;
				8'b1000101: c <= 9'b111001101;
				8'b1011001: c <= 9'b100000010;
				8'b110100: c <= 9'b110001100;
				8'b1111001: c <= 9'b101010000;
				8'b1110001: c <= 9'b10101000;
				8'b1001111: c <= 9'b10001010;
				8'b1100101: c <= 9'b111111000;
				8'b1111110: c <= 9'b10000101;
				8'b1111100: c <= 9'b10011101;
				8'b1010110: c <= 9'b11000110;
				8'b110010: c <= 9'b101110110;
				8'b1101101: c <= 9'b11101111;
				8'b100011: c <= 9'b11011101;
				8'b1110101: c <= 9'b100101111;
				8'b1111101: c <= 9'b111100101;
				8'b101001: c <= 9'b11001001;
				8'b1010010: c <= 9'b100111111;
				8'b1011000: c <= 9'b101110011;
				8'b101110: c <= 9'b111010110;
				8'b1000001: c <= 9'b10000111;
				default: c <= 9'b0;
			endcase
			9'b100000010 : case(di)
				8'b1000011: c <= 9'b11001;
				8'b101000: c <= 9'b11100111;
				8'b111010: c <= 9'b10011001;
				8'b110110: c <= 9'b110011011;
				8'b1100100: c <= 9'b11001111;
				8'b1000000: c <= 9'b110001110;
				8'b1110110: c <= 9'b111101010;
				8'b100101: c <= 9'b10100100;
				8'b101111: c <= 9'b100001100;
				8'b100110: c <= 9'b1111110;
				8'b1100011: c <= 9'b101100010;
				8'b1001000: c <= 9'b1101000;
				8'b111000: c <= 9'b1001101;
				8'b110001: c <= 9'b1110101;
				8'b1010111: c <= 9'b100111111;
				8'b1001110: c <= 9'b10100011;
				8'b1101010: c <= 9'b1000011;
				8'b1001001: c <= 9'b100100;
				8'b1100000: c <= 9'b10;
				8'b110111: c <= 9'b1000101;
				8'b1011101: c <= 9'b11000001;
				8'b1011011: c <= 9'b100111100;
				8'b111001: c <= 9'b10100110;
				8'b1001010: c <= 9'b11100010;
				8'b110011: c <= 9'b11111101;
				8'b1101100: c <= 9'b1001;
				8'b1110111: c <= 9'b10111110;
				8'b101011: c <= 9'b10000101;
				8'b1101011: c <= 9'b1001101;
				8'b111100: c <= 9'b110100101;
				8'b1000111: c <= 9'b101110111;
				8'b1011111: c <= 9'b11110011;
				8'b1110100: c <= 9'b100011111;
				8'b101101: c <= 9'b10000001;
				8'b1010011: c <= 9'b11001000;
				8'b1100001: c <= 9'b111010000;
				8'b110101: c <= 9'b1101111;
				8'b1000100: c <= 9'b110110;
				8'b1010001: c <= 9'b1010001;
				8'b1010100: c <= 9'b10011;
				8'b1100110: c <= 9'b10;
				8'b101010: c <= 9'b1111111;
				8'b1011110: c <= 9'b10111110;
				8'b1100111: c <= 9'b10110001;
				8'b1011010: c <= 9'b111101111;
				8'b1000010: c <= 9'b101100000;
				8'b111101: c <= 9'b110100110;
				8'b110000: c <= 9'b11011011;
				8'b111110: c <= 9'b10100000;
				8'b1100010: c <= 9'b100001001;
				8'b1110000: c <= 9'b100111000;
				8'b1101001: c <= 9'b100010011;
				8'b1110011: c <= 9'b101001110;
				8'b1001100: c <= 9'b10101011;
				8'b100001: c <= 9'b11010010;
				8'b1000110: c <= 9'b111110000;
				8'b1110010: c <= 9'b10011001;
				8'b1010000: c <= 9'b10011011;
				8'b1111010: c <= 9'b110101100;
				8'b1010101: c <= 9'b100001111;
				8'b111011: c <= 9'b1010011;
				8'b1001101: c <= 9'b1001011;
				8'b111111: c <= 9'b101101100;
				8'b1101110: c <= 9'b1101101;
				8'b1111011: c <= 9'b10001010;
				8'b1001011: c <= 9'b1000010;
				8'b1101111: c <= 9'b11011011;
				8'b1101000: c <= 9'b1111101;
				8'b101100: c <= 9'b1000111;
				8'b100100: c <= 9'b111100011;
				8'b1111000: c <= 9'b1110001;
				8'b1000101: c <= 9'b101001110;
				8'b1011001: c <= 9'b110101011;
				8'b110100: c <= 9'b1111010;
				8'b1111001: c <= 9'b10110011;
				8'b1110001: c <= 9'b11001111;
				8'b1001111: c <= 9'b110111111;
				8'b1100101: c <= 9'b110100;
				8'b1111110: c <= 9'b10010110;
				8'b1111100: c <= 9'b10010110;
				8'b1010110: c <= 9'b100000101;
				8'b110010: c <= 9'b1110001;
				8'b1101101: c <= 9'b110110011;
				8'b100011: c <= 9'b10000001;
				8'b1110101: c <= 9'b110110010;
				8'b1111101: c <= 9'b110110000;
				8'b101001: c <= 9'b11001110;
				8'b1010010: c <= 9'b111100;
				8'b1011000: c <= 9'b11010101;
				8'b101110: c <= 9'b100011010;
				8'b1000001: c <= 9'b11110111;
				default: c <= 9'b0;
			endcase
			9'b1111001 : case(di)
				8'b1000011: c <= 9'b111101010;
				8'b101000: c <= 9'b1110101;
				8'b111010: c <= 9'b11111000;
				8'b110110: c <= 9'b101001010;
				8'b1100100: c <= 9'b111111101;
				8'b1000000: c <= 9'b101110101;
				8'b1110110: c <= 9'b110100;
				8'b100101: c <= 9'b110000001;
				8'b101111: c <= 9'b1111101;
				8'b100110: c <= 9'b111001011;
				8'b1100011: c <= 9'b10111011;
				8'b1001000: c <= 9'b10011000;
				8'b111000: c <= 9'b111100111;
				8'b110001: c <= 9'b100101001;
				8'b1010111: c <= 9'b1100111;
				8'b1001110: c <= 9'b11100001;
				8'b1101010: c <= 9'b1010010;
				8'b1001001: c <= 9'b1100100;
				8'b1100000: c <= 9'b10101111;
				8'b110111: c <= 9'b1100010;
				8'b1011101: c <= 9'b100110101;
				8'b1011011: c <= 9'b11010;
				8'b111001: c <= 9'b10011010;
				8'b1001010: c <= 9'b100010;
				8'b110011: c <= 9'b11010010;
				8'b1101100: c <= 9'b110001000;
				8'b1110111: c <= 9'b110101001;
				8'b101011: c <= 9'b11011;
				8'b1101011: c <= 9'b1010010;
				8'b111100: c <= 9'b10000011;
				8'b1000111: c <= 9'b1001001;
				8'b1011111: c <= 9'b111000101;
				8'b1110100: c <= 9'b11011000;
				8'b101101: c <= 9'b110111111;
				8'b1010011: c <= 9'b111001100;
				8'b1100001: c <= 9'b10001000;
				8'b110101: c <= 9'b10100000;
				8'b1000100: c <= 9'b1000111;
				8'b1010001: c <= 9'b11010010;
				8'b1010100: c <= 9'b1000011;
				8'b1100110: c <= 9'b110000001;
				8'b101010: c <= 9'b111001111;
				8'b1011110: c <= 9'b101110;
				8'b1100111: c <= 9'b111100110;
				8'b1011010: c <= 9'b100100;
				8'b1000010: c <= 9'b100110000;
				8'b111101: c <= 9'b10110001;
				8'b110000: c <= 9'b100100001;
				8'b111110: c <= 9'b100010110;
				8'b1100010: c <= 9'b111101010;
				8'b1110000: c <= 9'b101011001;
				8'b1101001: c <= 9'b101110100;
				8'b1110011: c <= 9'b100000010;
				8'b1001100: c <= 9'b111101101;
				8'b100001: c <= 9'b110011111;
				8'b1000110: c <= 9'b110001111;
				8'b1110010: c <= 9'b1000111;
				8'b1010000: c <= 9'b10000111;
				8'b1111010: c <= 9'b110101010;
				8'b1010101: c <= 9'b10111011;
				8'b111011: c <= 9'b11110000;
				8'b1001101: c <= 9'b10110110;
				8'b111111: c <= 9'b100111011;
				8'b1101110: c <= 9'b101001011;
				8'b1111011: c <= 9'b111010110;
				8'b1001011: c <= 9'b10011101;
				8'b1101111: c <= 9'b10000000;
				8'b1101000: c <= 9'b10000001;
				8'b101100: c <= 9'b111010110;
				8'b100100: c <= 9'b11101100;
				8'b1111000: c <= 9'b100011101;
				8'b1000101: c <= 9'b11011001;
				8'b1011001: c <= 9'b100011011;
				8'b110100: c <= 9'b11011110;
				8'b1111001: c <= 9'b101010010;
				8'b1110001: c <= 9'b11110111;
				8'b1001111: c <= 9'b110111011;
				8'b1100101: c <= 9'b111101001;
				8'b1111110: c <= 9'b11011001;
				8'b1111100: c <= 9'b101100010;
				8'b1010110: c <= 9'b101011101;
				8'b110010: c <= 9'b111111011;
				8'b1101101: c <= 9'b110110111;
				8'b100011: c <= 9'b101000010;
				8'b1110101: c <= 9'b1110;
				8'b1111101: c <= 9'b100010101;
				8'b101001: c <= 9'b110110100;
				8'b1010010: c <= 9'b11111110;
				8'b1011000: c <= 9'b1101111;
				8'b101110: c <= 9'b11000100;
				8'b1000001: c <= 9'b1110001;
				default: c <= 9'b0;
			endcase
			9'b111010 : case(di)
				8'b1000011: c <= 9'b111001001;
				8'b101000: c <= 9'b110100;
				8'b111010: c <= 9'b11111001;
				8'b110110: c <= 9'b101101011;
				8'b1100100: c <= 9'b110100;
				8'b1000000: c <= 9'b101111110;
				8'b1110110: c <= 9'b100001100;
				8'b100101: c <= 9'b1000;
				8'b101111: c <= 9'b111011;
				8'b100110: c <= 9'b101011;
				8'b1100011: c <= 9'b100000011;
				8'b1001000: c <= 9'b11110111;
				8'b111000: c <= 9'b1110100;
				8'b110001: c <= 9'b110010111;
				8'b1010111: c <= 9'b111100100;
				8'b1001110: c <= 9'b11100101;
				8'b1101010: c <= 9'b1000;
				8'b1001001: c <= 9'b1100101;
				8'b1100000: c <= 9'b110110;
				8'b110111: c <= 9'b1010001;
				8'b1011101: c <= 9'b101001010;
				8'b1011011: c <= 9'b1111100;
				8'b111001: c <= 9'b110000001;
				8'b1001010: c <= 9'b11010000;
				8'b110011: c <= 9'b1110001;
				8'b1101100: c <= 9'b10001111;
				8'b1110111: c <= 9'b101101110;
				8'b101011: c <= 9'b110001111;
				8'b1101011: c <= 9'b100011001;
				8'b111100: c <= 9'b11101000;
				8'b1000111: c <= 9'b11010000;
				8'b1011111: c <= 9'b100100011;
				8'b1110100: c <= 9'b11110101;
				8'b101101: c <= 9'b11000;
				8'b1010011: c <= 9'b1110001;
				8'b1100001: c <= 9'b101110100;
				8'b110101: c <= 9'b110010;
				8'b1000100: c <= 9'b10101;
				8'b1010001: c <= 9'b100100101;
				8'b1010100: c <= 9'b11001100;
				8'b1100110: c <= 9'b100100101;
				8'b101010: c <= 9'b11100110;
				8'b1011110: c <= 9'b101011011;
				8'b1100111: c <= 9'b111010100;
				8'b1011010: c <= 9'b101101111;
				8'b1000010: c <= 9'b100011000;
				8'b111101: c <= 9'b10110100;
				8'b110000: c <= 9'b101101101;
				8'b111110: c <= 9'b110101100;
				8'b1100010: c <= 9'b10100010;
				8'b1110000: c <= 9'b10001111;
				8'b1101001: c <= 9'b11000000;
				8'b1110011: c <= 9'b1011010;
				8'b1001100: c <= 9'b11011011;
				8'b100001: c <= 9'b11001010;
				8'b1000110: c <= 9'b10011101;
				8'b1110010: c <= 9'b110000;
				8'b1010000: c <= 9'b111011101;
				8'b1111010: c <= 9'b1110011;
				8'b1010101: c <= 9'b111001100;
				8'b111011: c <= 9'b111010000;
				8'b1001101: c <= 9'b10110;
				8'b111111: c <= 9'b110100001;
				8'b1101110: c <= 9'b100001010;
				8'b1111011: c <= 9'b101110010;
				8'b1001011: c <= 9'b1000111;
				8'b1101111: c <= 9'b100110;
				8'b1101000: c <= 9'b101110011;
				8'b101100: c <= 9'b1100111;
				8'b100100: c <= 9'b1010011;
				8'b1111000: c <= 9'b10000;
				8'b1000101: c <= 9'b110101011;
				8'b1011001: c <= 9'b100111;
				8'b110100: c <= 9'b11010001;
				8'b1111001: c <= 9'b110000110;
				8'b1110001: c <= 9'b101001;
				8'b1001111: c <= 9'b101011111;
				8'b1100101: c <= 9'b11111;
				8'b1111110: c <= 9'b110000110;
				8'b1111100: c <= 9'b10110101;
				8'b1010110: c <= 9'b100101100;
				8'b110010: c <= 9'b100001110;
				8'b1101101: c <= 9'b100000001;
				8'b100011: c <= 9'b100010100;
				8'b1110101: c <= 9'b11010010;
				8'b1111101: c <= 9'b111110011;
				8'b101001: c <= 9'b11111000;
				8'b1010010: c <= 9'b110101100;
				8'b1011000: c <= 9'b10111001;
				8'b101110: c <= 9'b10001010;
				8'b1000001: c <= 9'b10000111;
				default: c <= 9'b0;
			endcase
			9'b110110010 : case(di)
				8'b1000011: c <= 9'b101010101;
				8'b101000: c <= 9'b101110001;
				8'b111010: c <= 9'b110010110;
				8'b110110: c <= 9'b1001111;
				8'b1100100: c <= 9'b11101;
				8'b1000000: c <= 9'b101001100;
				8'b1110110: c <= 9'b101000001;
				8'b100101: c <= 9'b1001010;
				8'b101111: c <= 9'b11101111;
				8'b100110: c <= 9'b111111111;
				8'b1100011: c <= 9'b11001100;
				8'b1001000: c <= 9'b110000110;
				8'b111000: c <= 9'b111000;
				8'b110001: c <= 9'b100110100;
				8'b1010111: c <= 9'b101100;
				8'b1001110: c <= 9'b111111001;
				8'b1101010: c <= 9'b1111011;
				8'b1001001: c <= 9'b101100;
				8'b1100000: c <= 9'b1110000;
				8'b110111: c <= 9'b1011011;
				8'b1011101: c <= 9'b10100;
				8'b1011011: c <= 9'b110110101;
				8'b111001: c <= 9'b11101100;
				8'b1001010: c <= 9'b101111000;
				8'b110011: c <= 9'b111001110;
				8'b1101100: c <= 9'b110010010;
				8'b1110111: c <= 9'b10000001;
				8'b101011: c <= 9'b110001010;
				8'b1101011: c <= 9'b100011;
				8'b111100: c <= 9'b1110;
				8'b1000111: c <= 9'b111011110;
				8'b1011111: c <= 9'b110101100;
				8'b1110100: c <= 9'b11010000;
				8'b101101: c <= 9'b11110001;
				8'b1010011: c <= 9'b11110000;
				8'b1100001: c <= 9'b10011001;
				8'b110101: c <= 9'b101000101;
				8'b1000100: c <= 9'b101;
				8'b1010001: c <= 9'b110011111;
				8'b1010100: c <= 9'b100011101;
				8'b1100110: c <= 9'b11101011;
				8'b101010: c <= 9'b11;
				8'b1011110: c <= 9'b1111000;
				8'b1100111: c <= 9'b111100010;
				8'b1011010: c <= 9'b110011000;
				8'b1000010: c <= 9'b100011000;
				8'b111101: c <= 9'b101100101;
				8'b110000: c <= 9'b100111010;
				8'b111110: c <= 9'b111101000;
				8'b1100010: c <= 9'b11100111;
				8'b1110000: c <= 9'b11101;
				8'b1101001: c <= 9'b111011011;
				8'b1110011: c <= 9'b110101010;
				8'b1001100: c <= 9'b100101010;
				8'b100001: c <= 9'b1110111;
				8'b1000110: c <= 9'b111001001;
				8'b1110010: c <= 9'b101011101;
				8'b1010000: c <= 9'b100000111;
				8'b1111010: c <= 9'b10101;
				8'b1010101: c <= 9'b10000111;
				8'b111011: c <= 9'b11011000;
				8'b1001101: c <= 9'b10110011;
				8'b111111: c <= 9'b111001001;
				8'b1101110: c <= 9'b111101111;
				8'b1111011: c <= 9'b11010000;
				8'b1001011: c <= 9'b100011010;
				8'b1101111: c <= 9'b110110000;
				8'b1101000: c <= 9'b110000110;
				8'b101100: c <= 9'b111101;
				8'b100100: c <= 9'b10111;
				8'b1111000: c <= 9'b100110000;
				8'b1000101: c <= 9'b10011000;
				8'b1011001: c <= 9'b110111110;
				8'b110100: c <= 9'b111000010;
				8'b1111001: c <= 9'b110111001;
				8'b1110001: c <= 9'b100010111;
				8'b1001111: c <= 9'b100001100;
				8'b1100101: c <= 9'b110101001;
				8'b1111110: c <= 9'b101110;
				8'b1111100: c <= 9'b1100;
				8'b1010110: c <= 9'b101010111;
				8'b110010: c <= 9'b11110100;
				8'b1101101: c <= 9'b10100111;
				8'b100011: c <= 9'b100111000;
				8'b1110101: c <= 9'b1111010;
				8'b1111101: c <= 9'b111110000;
				8'b101001: c <= 9'b100111110;
				8'b1010010: c <= 9'b111100000;
				8'b1011000: c <= 9'b111111001;
				8'b101110: c <= 9'b1000111;
				8'b1000001: c <= 9'b111001;
				default: c <= 9'b0;
			endcase
			9'b111001110 : case(di)
				8'b1000011: c <= 9'b110100111;
				8'b101000: c <= 9'b1000001;
				8'b111010: c <= 9'b110111000;
				8'b110110: c <= 9'b11100001;
				8'b1100100: c <= 9'b111010000;
				8'b1000000: c <= 9'b101001;
				8'b1110110: c <= 9'b100001110;
				8'b100101: c <= 9'b111010100;
				8'b101111: c <= 9'b101101;
				8'b100110: c <= 9'b110111010;
				8'b1100011: c <= 9'b1011000;
				8'b1001000: c <= 9'b111010100;
				8'b111000: c <= 9'b10000011;
				8'b110001: c <= 9'b1000000;
				8'b1010111: c <= 9'b110001;
				8'b1001110: c <= 9'b111101;
				8'b1101010: c <= 9'b100100011;
				8'b1001001: c <= 9'b110111000;
				8'b1100000: c <= 9'b111001110;
				8'b110111: c <= 9'b111000111;
				8'b1011101: c <= 9'b11101111;
				8'b1011011: c <= 9'b11101001;
				8'b111001: c <= 9'b100010101;
				8'b1001010: c <= 9'b101000110;
				8'b110011: c <= 9'b100001011;
				8'b1101100: c <= 9'b11001001;
				8'b1110111: c <= 9'b100101110;
				8'b101011: c <= 9'b101;
				8'b1101011: c <= 9'b11001000;
				8'b111100: c <= 9'b110001011;
				8'b1000111: c <= 9'b111000010;
				8'b1011111: c <= 9'b100000101;
				8'b1110100: c <= 9'b101001111;
				8'b101101: c <= 9'b110000010;
				8'b1010011: c <= 9'b1100011;
				8'b1100001: c <= 9'b11101101;
				8'b110101: c <= 9'b111010111;
				8'b1000100: c <= 9'b11001110;
				8'b1010001: c <= 9'b1000110;
				8'b1010100: c <= 9'b111101100;
				8'b1100110: c <= 9'b110101101;
				8'b101010: c <= 9'b100001010;
				8'b1011110: c <= 9'b11100000;
				8'b1100111: c <= 9'b11110111;
				8'b1011010: c <= 9'b110110;
				8'b1000010: c <= 9'b11000110;
				8'b111101: c <= 9'b11100001;
				8'b110000: c <= 9'b101001000;
				8'b111110: c <= 9'b101110;
				8'b1100010: c <= 9'b111000000;
				8'b1110000: c <= 9'b1101010;
				8'b1101001: c <= 9'b10111101;
				8'b1110011: c <= 9'b11000010;
				8'b1001100: c <= 9'b110000000;
				8'b100001: c <= 9'b111101110;
				8'b1000110: c <= 9'b10110;
				8'b1110010: c <= 9'b1111000;
				8'b1010000: c <= 9'b100111010;
				8'b1111010: c <= 9'b1101;
				8'b1010101: c <= 9'b10011100;
				8'b111011: c <= 9'b101101110;
				8'b1001101: c <= 9'b10101001;
				8'b111111: c <= 9'b111011101;
				8'b1101110: c <= 9'b101101010;
				8'b1111011: c <= 9'b110111;
				8'b1001011: c <= 9'b110010101;
				8'b1101111: c <= 9'b101001111;
				8'b1101000: c <= 9'b110110011;
				8'b101100: c <= 9'b11111010;
				8'b100100: c <= 9'b111011010;
				8'b1111000: c <= 9'b100010101;
				8'b1000101: c <= 9'b10010011;
				8'b1011001: c <= 9'b101101001;
				8'b110100: c <= 9'b10001110;
				8'b1111001: c <= 9'b11111000;
				8'b1110001: c <= 9'b110;
				8'b1001111: c <= 9'b1011010;
				8'b1100101: c <= 9'b110100111;
				8'b1111110: c <= 9'b110101111;
				8'b1111100: c <= 9'b11100110;
				8'b1010110: c <= 9'b101010100;
				8'b110010: c <= 9'b1101111;
				8'b1101101: c <= 9'b110010110;
				8'b100011: c <= 9'b10101111;
				8'b1110101: c <= 9'b1111110;
				8'b1111101: c <= 9'b100100010;
				8'b101001: c <= 9'b101010111;
				8'b1010010: c <= 9'b11010010;
				8'b1011000: c <= 9'b10011011;
				8'b101110: c <= 9'b100111010;
				8'b1000001: c <= 9'b10101101;
				default: c <= 9'b0;
			endcase
			9'b10011001 : case(di)
				8'b1000011: c <= 9'b110001011;
				8'b101000: c <= 9'b100111100;
				8'b111010: c <= 9'b11010001;
				8'b110110: c <= 9'b11010010;
				8'b1100100: c <= 9'b110100101;
				8'b1000000: c <= 9'b111110011;
				8'b1110110: c <= 9'b1100011;
				8'b100101: c <= 9'b10000111;
				8'b101111: c <= 9'b10111001;
				8'b100110: c <= 9'b10000011;
				8'b1100011: c <= 9'b111011010;
				8'b1001000: c <= 9'b100001010;
				8'b111000: c <= 9'b1110111;
				8'b110001: c <= 9'b101000010;
				8'b1010111: c <= 9'b10000011;
				8'b1001110: c <= 9'b10000;
				8'b1101010: c <= 9'b100110110;
				8'b1001001: c <= 9'b101101100;
				8'b1100000: c <= 9'b101110;
				8'b110111: c <= 9'b10000111;
				8'b1011101: c <= 9'b101110010;
				8'b1011011: c <= 9'b10111110;
				8'b111001: c <= 9'b10110;
				8'b1001010: c <= 9'b101100100;
				8'b110011: c <= 9'b11000100;
				8'b1101100: c <= 9'b1101111;
				8'b1110111: c <= 9'b100101000;
				8'b101011: c <= 9'b1001101;
				8'b1101011: c <= 9'b111000011;
				8'b111100: c <= 9'b10101000;
				8'b1000111: c <= 9'b1110000;
				8'b1011111: c <= 9'b111001101;
				8'b1110100: c <= 9'b111001110;
				8'b101101: c <= 9'b100000100;
				8'b1010011: c <= 9'b1011011;
				8'b1100001: c <= 9'b101010011;
				8'b110101: c <= 9'b101011110;
				8'b1000100: c <= 9'b111010110;
				8'b1010001: c <= 9'b11010001;
				8'b1010100: c <= 9'b11011001;
				8'b1100110: c <= 9'b111000000;
				8'b101010: c <= 9'b101000011;
				8'b1011110: c <= 9'b111010001;
				8'b1100111: c <= 9'b110000101;
				8'b1011010: c <= 9'b1000000;
				8'b1000010: c <= 9'b101101001;
				8'b111101: c <= 9'b111100110;
				8'b110000: c <= 9'b11101011;
				8'b111110: c <= 9'b100010;
				8'b1100010: c <= 9'b1110100;
				8'b1110000: c <= 9'b10010011;
				8'b1101001: c <= 9'b100010010;
				8'b1110011: c <= 9'b11010011;
				8'b1001100: c <= 9'b10111000;
				8'b100001: c <= 9'b11110001;
				8'b1000110: c <= 9'b1110010;
				8'b1110010: c <= 9'b1100110;
				8'b1010000: c <= 9'b11111010;
				8'b1111010: c <= 9'b101001000;
				8'b1010101: c <= 9'b101010010;
				8'b111011: c <= 9'b1000011;
				8'b1001101: c <= 9'b111010;
				8'b111111: c <= 9'b110011100;
				8'b1101110: c <= 9'b10101000;
				8'b1111011: c <= 9'b111111101;
				8'b1001011: c <= 9'b111001000;
				8'b1101111: c <= 9'b11100111;
				8'b1101000: c <= 9'b110001000;
				8'b101100: c <= 9'b100010000;
				8'b100100: c <= 9'b100100;
				8'b1111000: c <= 9'b101001010;
				8'b1000101: c <= 9'b101111010;
				8'b1011001: c <= 9'b111100100;
				8'b110100: c <= 9'b110101101;
				8'b1111001: c <= 9'b10011100;
				8'b1110001: c <= 9'b110011001;
				8'b1001111: c <= 9'b10010110;
				8'b1100101: c <= 9'b111111110;
				8'b1111110: c <= 9'b100011011;
				8'b1111100: c <= 9'b110110010;
				8'b1010110: c <= 9'b1101110;
				8'b110010: c <= 9'b101110111;
				8'b1101101: c <= 9'b110000111;
				8'b100011: c <= 9'b1001101;
				8'b1110101: c <= 9'b100101100;
				8'b1111101: c <= 9'b110011001;
				8'b101001: c <= 9'b10011100;
				8'b1010010: c <= 9'b10000111;
				8'b1011000: c <= 9'b100101100;
				8'b101110: c <= 9'b10010000;
				8'b1000001: c <= 9'b11100100;
				default: c <= 9'b0;
			endcase
			9'b101010100 : case(di)
				8'b1000011: c <= 9'b101000010;
				8'b101000: c <= 9'b1110001;
				8'b111010: c <= 9'b1111011;
				8'b110110: c <= 9'b1000;
				8'b1100100: c <= 9'b1100;
				8'b1000000: c <= 9'b101001111;
				8'b1110110: c <= 9'b10101110;
				8'b100101: c <= 9'b101111001;
				8'b101111: c <= 9'b111101010;
				8'b100110: c <= 9'b101000010;
				8'b1100011: c <= 9'b101000011;
				8'b1001000: c <= 9'b111101;
				8'b111000: c <= 9'b110100111;
				8'b110001: c <= 9'b111111110;
				8'b1010111: c <= 9'b10101100;
				8'b1001110: c <= 9'b1111000;
				8'b1101010: c <= 9'b110100;
				8'b1001001: c <= 9'b110000001;
				8'b1100000: c <= 9'b1011000;
				8'b110111: c <= 9'b100111000;
				8'b1011101: c <= 9'b101001010;
				8'b1011011: c <= 9'b100000000;
				8'b111001: c <= 9'b110100111;
				8'b1001010: c <= 9'b111010;
				8'b110011: c <= 9'b100110100;
				8'b1101100: c <= 9'b100001;
				8'b1110111: c <= 9'b111010110;
				8'b101011: c <= 9'b11011001;
				8'b1101011: c <= 9'b110111011;
				8'b111100: c <= 9'b101101;
				8'b1000111: c <= 9'b110110000;
				8'b1011111: c <= 9'b101001110;
				8'b1110100: c <= 9'b10000111;
				8'b101101: c <= 9'b100101100;
				8'b1010011: c <= 9'b110000001;
				8'b1100001: c <= 9'b100011100;
				8'b110101: c <= 9'b101001011;
				8'b1000100: c <= 9'b100010000;
				8'b1010001: c <= 9'b111011101;
				8'b1010100: c <= 9'b10100011;
				8'b1100110: c <= 9'b101101011;
				8'b101010: c <= 9'b1100101;
				8'b1011110: c <= 9'b111011101;
				8'b1100111: c <= 9'b110011111;
				8'b1011010: c <= 9'b101111000;
				8'b1000010: c <= 9'b111011010;
				8'b111101: c <= 9'b11101011;
				8'b110000: c <= 9'b100111111;
				8'b111110: c <= 9'b100010000;
				8'b1100010: c <= 9'b10011010;
				8'b1110000: c <= 9'b10;
				8'b1101001: c <= 9'b101101101;
				8'b1110011: c <= 9'b111001;
				8'b1001100: c <= 9'b101101100;
				8'b100001: c <= 9'b111110101;
				8'b1000110: c <= 9'b11001110;
				8'b1110010: c <= 9'b11111000;
				8'b1010000: c <= 9'b10110010;
				8'b1111010: c <= 9'b11001100;
				8'b1010101: c <= 9'b100011101;
				8'b111011: c <= 9'b101101010;
				8'b1001101: c <= 9'b10011000;
				8'b111111: c <= 9'b101110100;
				8'b1101110: c <= 9'b1110011;
				8'b1111011: c <= 9'b100110111;
				8'b1001011: c <= 9'b100010010;
				8'b1101111: c <= 9'b1111010;
				8'b1101000: c <= 9'b100110111;
				8'b101100: c <= 9'b100;
				8'b100100: c <= 9'b100010011;
				8'b1111000: c <= 9'b1111111;
				8'b1000101: c <= 9'b101101000;
				8'b1011001: c <= 9'b10001011;
				8'b110100: c <= 9'b101110101;
				8'b1111001: c <= 9'b110000111;
				8'b1110001: c <= 9'b110101111;
				8'b1001111: c <= 9'b10101111;
				8'b1100101: c <= 9'b10010110;
				8'b1111110: c <= 9'b11001001;
				8'b1111100: c <= 9'b101101;
				8'b1010110: c <= 9'b11011000;
				8'b110010: c <= 9'b10110001;
				8'b1101101: c <= 9'b110010100;
				8'b100011: c <= 9'b10101000;
				8'b1110101: c <= 9'b100100111;
				8'b1111101: c <= 9'b10100110;
				8'b101001: c <= 9'b110011011;
				8'b1010010: c <= 9'b111011100;
				8'b1011000: c <= 9'b100000001;
				8'b101110: c <= 9'b11100101;
				8'b1000001: c <= 9'b11100100;
				default: c <= 9'b0;
			endcase
			9'b10111010 : case(di)
				8'b1000011: c <= 9'b10000011;
				8'b101000: c <= 9'b1101010;
				8'b111010: c <= 9'b110011010;
				8'b110110: c <= 9'b101000001;
				8'b1100100: c <= 9'b110100001;
				8'b1000000: c <= 9'b101001110;
				8'b1110110: c <= 9'b110001010;
				8'b100101: c <= 9'b1000;
				8'b101111: c <= 9'b101100;
				8'b100110: c <= 9'b110100010;
				8'b1100011: c <= 9'b111100110;
				8'b1001000: c <= 9'b110011010;
				8'b111000: c <= 9'b101111000;
				8'b110001: c <= 9'b111011010;
				8'b1010111: c <= 9'b11111001;
				8'b1001110: c <= 9'b100010000;
				8'b1101010: c <= 9'b10100101;
				8'b1001001: c <= 9'b10010011;
				8'b1100000: c <= 9'b110000010;
				8'b110111: c <= 9'b100010101;
				8'b1011101: c <= 9'b11011101;
				8'b1011011: c <= 9'b110110100;
				8'b111001: c <= 9'b101110101;
				8'b1001010: c <= 9'b101011000;
				8'b110011: c <= 9'b110101;
				8'b1101100: c <= 9'b110000110;
				8'b1110111: c <= 9'b111010010;
				8'b101011: c <= 9'b10100101;
				8'b1101011: c <= 9'b101110010;
				8'b111100: c <= 9'b10000111;
				8'b1000111: c <= 9'b100000010;
				8'b1011111: c <= 9'b10111100;
				8'b1110100: c <= 9'b110;
				8'b101101: c <= 9'b110111010;
				8'b1010011: c <= 9'b111111011;
				8'b1100001: c <= 9'b100110110;
				8'b110101: c <= 9'b11101000;
				8'b1000100: c <= 9'b11111100;
				8'b1010001: c <= 9'b110110100;
				8'b1010100: c <= 9'b100000000;
				8'b1100110: c <= 9'b1100011;
				8'b101010: c <= 9'b11110110;
				8'b1011110: c <= 9'b111101110;
				8'b1100111: c <= 9'b110100111;
				8'b1011010: c <= 9'b1001101;
				8'b1000010: c <= 9'b111101000;
				8'b111101: c <= 9'b1001010;
				8'b110000: c <= 9'b11100111;
				8'b111110: c <= 9'b100111010;
				8'b1100010: c <= 9'b111000;
				8'b1110000: c <= 9'b100111011;
				8'b1101001: c <= 9'b111001111;
				8'b1110011: c <= 9'b100001010;
				8'b1001100: c <= 9'b111010100;
				8'b100001: c <= 9'b101100101;
				8'b1000110: c <= 9'b10000111;
				8'b1110010: c <= 9'b110001110;
				8'b1010000: c <= 9'b101011111;
				8'b1111010: c <= 9'b110010101;
				8'b1010101: c <= 9'b110110;
				8'b111011: c <= 9'b11110111;
				8'b1001101: c <= 9'b110011100;
				8'b111111: c <= 9'b11010001;
				8'b1101110: c <= 9'b10000011;
				8'b1111011: c <= 9'b1101101;
				8'b1001011: c <= 9'b1011111;
				8'b1101111: c <= 9'b111100100;
				8'b1101000: c <= 9'b101111010;
				8'b101100: c <= 9'b10110110;
				8'b100100: c <= 9'b101001100;
				8'b1111000: c <= 9'b110100011;
				8'b1000101: c <= 9'b10101011;
				8'b1011001: c <= 9'b1111100;
				8'b110100: c <= 9'b11111011;
				8'b1111001: c <= 9'b101110100;
				8'b1110001: c <= 9'b100010111;
				8'b1001111: c <= 9'b111000101;
				8'b1100101: c <= 9'b11110;
				8'b1111110: c <= 9'b111100000;
				8'b1111100: c <= 9'b111001101;
				8'b1010110: c <= 9'b111101001;
				8'b110010: c <= 9'b110101110;
				8'b1101101: c <= 9'b11110001;
				8'b100011: c <= 9'b100110;
				8'b1110101: c <= 9'b10010110;
				8'b1111101: c <= 9'b100001101;
				8'b101001: c <= 9'b101010000;
				8'b1010010: c <= 9'b1111110;
				8'b1011000: c <= 9'b100001011;
				8'b101110: c <= 9'b101011001;
				8'b1000001: c <= 9'b100100;
				default: c <= 9'b0;
			endcase
			9'b11011110 : case(di)
				8'b1000011: c <= 9'b110110000;
				8'b101000: c <= 9'b110011101;
				8'b111010: c <= 9'b110111010;
				8'b110110: c <= 9'b101000110;
				8'b1100100: c <= 9'b11111010;
				8'b1000000: c <= 9'b110010100;
				8'b1110110: c <= 9'b11100011;
				8'b100101: c <= 9'b10010;
				8'b101111: c <= 9'b110000;
				8'b100110: c <= 9'b11010011;
				8'b1100011: c <= 9'b10100111;
				8'b1001000: c <= 9'b10010111;
				8'b111000: c <= 9'b111001111;
				8'b110001: c <= 9'b100100101;
				8'b1010111: c <= 9'b1100010;
				8'b1001110: c <= 9'b11011010;
				8'b1101010: c <= 9'b111101001;
				8'b1001001: c <= 9'b1010110;
				8'b1100000: c <= 9'b10001011;
				8'b110111: c <= 9'b11001000;
				8'b1011101: c <= 9'b100010101;
				8'b1011011: c <= 9'b110010001;
				8'b111001: c <= 9'b110110100;
				8'b1001010: c <= 9'b10010101;
				8'b110011: c <= 9'b1110111;
				8'b1101100: c <= 9'b101101110;
				8'b1110111: c <= 9'b110111011;
				8'b101011: c <= 9'b10011111;
				8'b1101011: c <= 9'b100110011;
				8'b111100: c <= 9'b111011011;
				8'b1000111: c <= 9'b110000;
				8'b1011111: c <= 9'b11000;
				8'b1110100: c <= 9'b101100101;
				8'b101101: c <= 9'b11001;
				8'b1010011: c <= 9'b111000100;
				8'b1100001: c <= 9'b101001100;
				8'b110101: c <= 9'b111011010;
				8'b1000100: c <= 9'b1100100;
				8'b1010001: c <= 9'b100110100;
				8'b1010100: c <= 9'b101100100;
				8'b1100110: c <= 9'b101011111;
				8'b101010: c <= 9'b100100011;
				8'b1011110: c <= 9'b100110;
				8'b1100111: c <= 9'b11001011;
				8'b1011010: c <= 9'b1001110;
				8'b1000010: c <= 9'b11000111;
				8'b111101: c <= 9'b100111100;
				8'b110000: c <= 9'b110100;
				8'b111110: c <= 9'b101100010;
				8'b1100010: c <= 9'b10100101;
				8'b1110000: c <= 9'b101101111;
				8'b1101001: c <= 9'b111000000;
				8'b1110011: c <= 9'b110001101;
				8'b1001100: c <= 9'b110110;
				8'b100001: c <= 9'b111000011;
				8'b1000110: c <= 9'b11000;
				8'b1110010: c <= 9'b111110110;
				8'b1010000: c <= 9'b110001;
				8'b1111010: c <= 9'b100101001;
				8'b1010101: c <= 9'b100111000;
				8'b111011: c <= 9'b11001011;
				8'b1001101: c <= 9'b10010100;
				8'b111111: c <= 9'b10011010;
				8'b1101110: c <= 9'b10111;
				8'b1111011: c <= 9'b100100;
				8'b1001011: c <= 9'b111000100;
				8'b1101111: c <= 9'b10111110;
				8'b1101000: c <= 9'b110000110;
				8'b101100: c <= 9'b111101110;
				8'b100100: c <= 9'b101111010;
				8'b1111000: c <= 9'b101101111;
				8'b1000101: c <= 9'b100100;
				8'b1011001: c <= 9'b100101000;
				8'b110100: c <= 9'b1100;
				8'b1111001: c <= 9'b100111;
				8'b1110001: c <= 9'b10001110;
				8'b1001111: c <= 9'b111010100;
				8'b1100101: c <= 9'b1000111;
				8'b1111110: c <= 9'b111111111;
				8'b1111100: c <= 9'b110010;
				8'b1010110: c <= 9'b10101110;
				8'b110010: c <= 9'b10010111;
				8'b1101101: c <= 9'b101000011;
				8'b100011: c <= 9'b100101001;
				8'b1110101: c <= 9'b100010010;
				8'b1111101: c <= 9'b10010101;
				8'b101001: c <= 9'b110000000;
				8'b1010010: c <= 9'b100100101;
				8'b1011000: c <= 9'b110011111;
				8'b101110: c <= 9'b101000011;
				8'b1000001: c <= 9'b11111011;
				default: c <= 9'b0;
			endcase
			9'b111000110 : case(di)
				8'b1000011: c <= 9'b110101010;
				8'b101000: c <= 9'b101110;
				8'b111010: c <= 9'b11101001;
				8'b110110: c <= 9'b101001000;
				8'b1100100: c <= 9'b110110110;
				8'b1000000: c <= 9'b11110011;
				8'b1110110: c <= 9'b10111000;
				8'b100101: c <= 9'b10000011;
				8'b101111: c <= 9'b111001111;
				8'b100110: c <= 9'b11100;
				8'b1100011: c <= 9'b11000110;
				8'b1001000: c <= 9'b110101110;
				8'b111000: c <= 9'b1001110;
				8'b110001: c <= 9'b110110100;
				8'b1010111: c <= 9'b1001100;
				8'b1001110: c <= 9'b111010100;
				8'b1101010: c <= 9'b10100110;
				8'b1001001: c <= 9'b10011;
				8'b1100000: c <= 9'b11101001;
				8'b110111: c <= 9'b11100111;
				8'b1011101: c <= 9'b10111001;
				8'b1011011: c <= 9'b10100011;
				8'b111001: c <= 9'b111000101;
				8'b1001010: c <= 9'b10111011;
				8'b110011: c <= 9'b110110000;
				8'b1101100: c <= 9'b101101110;
				8'b1110111: c <= 9'b111010001;
				8'b101011: c <= 9'b101001010;
				8'b1101011: c <= 9'b100;
				8'b111100: c <= 9'b100010001;
				8'b1000111: c <= 9'b111010;
				8'b1011111: c <= 9'b10110010;
				8'b1110100: c <= 9'b100100001;
				8'b101101: c <= 9'b110010;
				8'b1010011: c <= 9'b10010011;
				8'b1100001: c <= 9'b100100000;
				8'b110101: c <= 9'b11100000;
				8'b1000100: c <= 9'b10110011;
				8'b1010001: c <= 9'b1110;
				8'b1010100: c <= 9'b10000010;
				8'b1100110: c <= 9'b110111010;
				8'b101010: c <= 9'b100111101;
				8'b1011110: c <= 9'b1000000;
				8'b1100111: c <= 9'b100110000;
				8'b1011010: c <= 9'b100111101;
				8'b1000010: c <= 9'b10001010;
				8'b111101: c <= 9'b110100100;
				8'b110000: c <= 9'b1111110;
				8'b111110: c <= 9'b1000;
				8'b1100010: c <= 9'b100001;
				8'b1110000: c <= 9'b111;
				8'b1101001: c <= 9'b11011001;
				8'b1110011: c <= 9'b110000000;
				8'b1001100: c <= 9'b110101100;
				8'b100001: c <= 9'b1000100;
				8'b1000110: c <= 9'b11111110;
				8'b1110010: c <= 9'b11001110;
				8'b1010000: c <= 9'b1111;
				8'b1111010: c <= 9'b11110010;
				8'b1010101: c <= 9'b1001000;
				8'b111011: c <= 9'b101101011;
				8'b1001101: c <= 9'b100110110;
				8'b111111: c <= 9'b110010100;
				8'b1101110: c <= 9'b11001;
				8'b1111011: c <= 9'b10101101;
				8'b1001011: c <= 9'b111101100;
				8'b1101111: c <= 9'b111000101;
				8'b1101000: c <= 9'b111111001;
				8'b101100: c <= 9'b110011011;
				8'b100100: c <= 9'b111011110;
				8'b1111000: c <= 9'b111000;
				8'b1000101: c <= 9'b101010001;
				8'b1011001: c <= 9'b11;
				8'b110100: c <= 9'b111111011;
				8'b1111001: c <= 9'b100110011;
				8'b1110001: c <= 9'b100101101;
				8'b1001111: c <= 9'b110011011;
				8'b1100101: c <= 9'b1101000;
				8'b1111110: c <= 9'b11100101;
				8'b1111100: c <= 9'b10011;
				8'b1010110: c <= 9'b111111011;
				8'b110010: c <= 9'b111100100;
				8'b1101101: c <= 9'b101000011;
				8'b100011: c <= 9'b11110000;
				8'b1110101: c <= 9'b101000;
				8'b1111101: c <= 9'b11010001;
				8'b101001: c <= 9'b110100011;
				8'b1010010: c <= 9'b10011100;
				8'b1011000: c <= 9'b111101110;
				8'b101110: c <= 9'b101101011;
				8'b1000001: c <= 9'b1111101;
				default: c <= 9'b0;
			endcase
			9'b10011011 : case(di)
				8'b1000011: c <= 9'b1111110;
				8'b101000: c <= 9'b100001010;
				8'b111010: c <= 9'b11010010;
				8'b110110: c <= 9'b11010111;
				8'b1100100: c <= 9'b1111011;
				8'b1000000: c <= 9'b111011101;
				8'b1110110: c <= 9'b11100000;
				8'b100101: c <= 9'b10001011;
				8'b101111: c <= 9'b101100010;
				8'b100110: c <= 9'b101000010;
				8'b1100011: c <= 9'b10010011;
				8'b1001000: c <= 9'b110100111;
				8'b111000: c <= 9'b1011010;
				8'b110001: c <= 9'b1000101;
				8'b1010111: c <= 9'b10001010;
				8'b1001110: c <= 9'b101100110;
				8'b1101010: c <= 9'b10101101;
				8'b1001001: c <= 9'b10001011;
				8'b1100000: c <= 9'b10010100;
				8'b110111: c <= 9'b10110011;
				8'b1011101: c <= 9'b110011111;
				8'b1011011: c <= 9'b111011111;
				8'b111001: c <= 9'b101110111;
				8'b1001010: c <= 9'b110011000;
				8'b110011: c <= 9'b1000;
				8'b1101100: c <= 9'b100011001;
				8'b1110111: c <= 9'b100110111;
				8'b101011: c <= 9'b101000100;
				8'b1101011: c <= 9'b101110001;
				8'b111100: c <= 9'b10100000;
				8'b1000111: c <= 9'b100010111;
				8'b1011111: c <= 9'b111101111;
				8'b1110100: c <= 9'b10100110;
				8'b101101: c <= 9'b1000110;
				8'b1010011: c <= 9'b110010011;
				8'b1100001: c <= 9'b101000110;
				8'b110101: c <= 9'b110101101;
				8'b1000100: c <= 9'b101010;
				8'b1010001: c <= 9'b1110101;
				8'b1010100: c <= 9'b10110100;
				8'b1100110: c <= 9'b100111100;
				8'b101010: c <= 9'b100000000;
				8'b1011110: c <= 9'b100100;
				8'b1100111: c <= 9'b100001010;
				8'b1011010: c <= 9'b101100101;
				8'b1000010: c <= 9'b101011;
				8'b111101: c <= 9'b100001001;
				8'b110000: c <= 9'b110100110;
				8'b111110: c <= 9'b101010101;
				8'b1100010: c <= 9'b1001101;
				8'b1110000: c <= 9'b111111111;
				8'b1101001: c <= 9'b1100;
				8'b1110011: c <= 9'b1111101;
				8'b1001100: c <= 9'b101010111;
				8'b100001: c <= 9'b110110111;
				8'b1000110: c <= 9'b101110000;
				8'b1110010: c <= 9'b100111100;
				8'b1010000: c <= 9'b111011011;
				8'b1111010: c <= 9'b10011111;
				8'b1010101: c <= 9'b1100011;
				8'b111011: c <= 9'b10101110;
				8'b1001101: c <= 9'b110010111;
				8'b111111: c <= 9'b11000001;
				8'b1101110: c <= 9'b110110110;
				8'b1111011: c <= 9'b11111101;
				8'b1001011: c <= 9'b1010101;
				8'b1101111: c <= 9'b1111011;
				8'b1101000: c <= 9'b1111011;
				8'b101100: c <= 9'b10110101;
				8'b100100: c <= 9'b10011000;
				8'b1111000: c <= 9'b101101111;
				8'b1000101: c <= 9'b110101001;
				8'b1011001: c <= 9'b1001101;
				8'b110100: c <= 9'b111100;
				8'b1111001: c <= 9'b101010000;
				8'b1110001: c <= 9'b10010;
				8'b1001111: c <= 9'b1100010;
				8'b1100101: c <= 9'b11100000;
				8'b1111110: c <= 9'b101010;
				8'b1111100: c <= 9'b110010111;
				8'b1010110: c <= 9'b111111010;
				8'b110010: c <= 9'b1111000;
				8'b1101101: c <= 9'b1001110;
				8'b100011: c <= 9'b100100;
				8'b1110101: c <= 9'b101000001;
				8'b1111101: c <= 9'b11100;
				8'b101001: c <= 9'b100110110;
				8'b1010010: c <= 9'b10000111;
				8'b1011000: c <= 9'b1010001;
				8'b101110: c <= 9'b111101001;
				8'b1000001: c <= 9'b11000001;
				default: c <= 9'b0;
			endcase
			9'b110100101 : case(di)
				8'b1000011: c <= 9'b100111100;
				8'b101000: c <= 9'b111110000;
				8'b111010: c <= 9'b10110001;
				8'b110110: c <= 9'b100000100;
				8'b1100100: c <= 9'b101110101;
				8'b1000000: c <= 9'b10000011;
				8'b1110110: c <= 9'b10111000;
				8'b100101: c <= 9'b110110110;
				8'b101111: c <= 9'b111000100;
				8'b100110: c <= 9'b100100;
				8'b1100011: c <= 9'b1001101;
				8'b1001000: c <= 9'b1100111;
				8'b111000: c <= 9'b1011;
				8'b110001: c <= 9'b10110101;
				8'b1010111: c <= 9'b1010011;
				8'b1001110: c <= 9'b1110001;
				8'b1101010: c <= 9'b1010101;
				8'b1001001: c <= 9'b1101;
				8'b1100000: c <= 9'b110010001;
				8'b110111: c <= 9'b111111110;
				8'b1011101: c <= 9'b10011001;
				8'b1011011: c <= 9'b111101;
				8'b111001: c <= 9'b10110110;
				8'b1001010: c <= 9'b10100111;
				8'b110011: c <= 9'b110000001;
				8'b1101100: c <= 9'b100100001;
				8'b1110111: c <= 9'b10111001;
				8'b101011: c <= 9'b1101;
				8'b1101011: c <= 9'b100111000;
				8'b111100: c <= 9'b1011111;
				8'b1000111: c <= 9'b101110001;
				8'b1011111: c <= 9'b101101011;
				8'b1110100: c <= 9'b1000100;
				8'b101101: c <= 9'b11100110;
				8'b1010011: c <= 9'b1101;
				8'b1100001: c <= 9'b110010010;
				8'b110101: c <= 9'b1111101;
				8'b1000100: c <= 9'b10100101;
				8'b1010001: c <= 9'b11101000;
				8'b1010100: c <= 9'b100;
				8'b1100110: c <= 9'b100100000;
				8'b101010: c <= 9'b10100011;
				8'b1011110: c <= 9'b10010100;
				8'b1100111: c <= 9'b101000100;
				8'b1011010: c <= 9'b11100110;
				8'b1000010: c <= 9'b10000110;
				8'b111101: c <= 9'b11001000;
				8'b110000: c <= 9'b10010100;
				8'b111110: c <= 9'b111101;
				8'b1100010: c <= 9'b101011101;
				8'b1110000: c <= 9'b111001001;
				8'b1101001: c <= 9'b1001011;
				8'b1110011: c <= 9'b111000000;
				8'b1001100: c <= 9'b10110110;
				8'b100001: c <= 9'b100001110;
				8'b1000110: c <= 9'b110010011;
				8'b1110010: c <= 9'b111110110;
				8'b1010000: c <= 9'b111000111;
				8'b1111010: c <= 9'b1110010;
				8'b1010101: c <= 9'b100000101;
				8'b111011: c <= 9'b100111100;
				8'b1001101: c <= 9'b11010001;
				8'b111111: c <= 9'b111001001;
				8'b1101110: c <= 9'b11010001;
				8'b1111011: c <= 9'b111101100;
				8'b1001011: c <= 9'b111010110;
				8'b1101111: c <= 9'b110;
				8'b1101000: c <= 9'b10100111;
				8'b101100: c <= 9'b11111001;
				8'b100100: c <= 9'b10100111;
				8'b1111000: c <= 9'b110111011;
				8'b1000101: c <= 9'b1110011;
				8'b1011001: c <= 9'b110011010;
				8'b110100: c <= 9'b111000101;
				8'b1111001: c <= 9'b110100110;
				8'b1110001: c <= 9'b11100101;
				8'b1001111: c <= 9'b11100110;
				8'b1100101: c <= 9'b111111111;
				8'b1111110: c <= 9'b100011111;
				8'b1111100: c <= 9'b10111000;
				8'b1010110: c <= 9'b110010110;
				8'b110010: c <= 9'b1000;
				8'b1101101: c <= 9'b11100010;
				8'b100011: c <= 9'b1110011;
				8'b1110101: c <= 9'b101011010;
				8'b1111101: c <= 9'b11110101;
				8'b101001: c <= 9'b111111111;
				8'b1010010: c <= 9'b11101100;
				8'b1011000: c <= 9'b1001110;
				8'b101110: c <= 9'b110001010;
				8'b1000001: c <= 9'b110100000;
				default: c <= 9'b0;
			endcase
			9'b110000010 : case(di)
				8'b1000011: c <= 9'b101000101;
				8'b101000: c <= 9'b100101111;
				8'b111010: c <= 9'b11011001;
				8'b110110: c <= 9'b101100111;
				8'b1100100: c <= 9'b101010;
				8'b1000000: c <= 9'b1001010;
				8'b1110110: c <= 9'b111101110;
				8'b100101: c <= 9'b10000000;
				8'b101111: c <= 9'b10110001;
				8'b100110: c <= 9'b100110100;
				8'b1100011: c <= 9'b101110000;
				8'b1001000: c <= 9'b11111010;
				8'b111000: c <= 9'b10000001;
				8'b110001: c <= 9'b100010010;
				8'b1010111: c <= 9'b11010;
				8'b1001110: c <= 9'b100101111;
				8'b1101010: c <= 9'b1011010;
				8'b1001001: c <= 9'b1100;
				8'b1100000: c <= 9'b101110100;
				8'b110111: c <= 9'b110111001;
				8'b1011101: c <= 9'b110011101;
				8'b1011011: c <= 9'b10111010;
				8'b111001: c <= 9'b100000110;
				8'b1001010: c <= 9'b110011101;
				8'b110011: c <= 9'b11010001;
				8'b1101100: c <= 9'b110000;
				8'b1110111: c <= 9'b111011110;
				8'b101011: c <= 9'b1101000;
				8'b1101011: c <= 9'b10001011;
				8'b111100: c <= 9'b110011010;
				8'b1000111: c <= 9'b10000101;
				8'b1011111: c <= 9'b100010000;
				8'b1110100: c <= 9'b101001;
				8'b101101: c <= 9'b101110010;
				8'b1010011: c <= 9'b10111001;
				8'b1100001: c <= 9'b10110001;
				8'b110101: c <= 9'b11000010;
				8'b1000100: c <= 9'b11010000;
				8'b1010001: c <= 9'b10100011;
				8'b1010100: c <= 9'b111100101;
				8'b1100110: c <= 9'b11011100;
				8'b101010: c <= 9'b10010111;
				8'b1011110: c <= 9'b100000010;
				8'b1100111: c <= 9'b101000101;
				8'b1011010: c <= 9'b10110011;
				8'b1000010: c <= 9'b101000101;
				8'b111101: c <= 9'b110000110;
				8'b110000: c <= 9'b1111010;
				8'b111110: c <= 9'b110101;
				8'b1100010: c <= 9'b110100101;
				8'b1110000: c <= 9'b101101110;
				8'b1101001: c <= 9'b100011100;
				8'b1110011: c <= 9'b10111000;
				8'b1001100: c <= 9'b11111110;
				8'b100001: c <= 9'b101101101;
				8'b1000110: c <= 9'b110001101;
				8'b1110010: c <= 9'b111001111;
				8'b1010000: c <= 9'b100100110;
				8'b1111010: c <= 9'b111001110;
				8'b1010101: c <= 9'b110111001;
				8'b111011: c <= 9'b11001001;
				8'b1001101: c <= 9'b10111000;
				8'b111111: c <= 9'b100011111;
				8'b1101110: c <= 9'b111001001;
				8'b1111011: c <= 9'b10001101;
				8'b1001011: c <= 9'b1010000;
				8'b1101111: c <= 9'b110000111;
				8'b1101000: c <= 9'b101110111;
				8'b101100: c <= 9'b10000101;
				8'b100100: c <= 9'b110101011;
				8'b1111000: c <= 9'b111011001;
				8'b1000101: c <= 9'b1010001;
				8'b1011001: c <= 9'b10100;
				8'b110100: c <= 9'b10010110;
				8'b1111001: c <= 9'b11101011;
				8'b1110001: c <= 9'b101111111;
				8'b1001111: c <= 9'b110011111;
				8'b1100101: c <= 9'b10111101;
				8'b1111110: c <= 9'b10101010;
				8'b1111100: c <= 9'b10110011;
				8'b1010110: c <= 9'b100110011;
				8'b110010: c <= 9'b11010100;
				8'b1101101: c <= 9'b100011;
				8'b100011: c <= 9'b11111101;
				8'b1110101: c <= 9'b101101101;
				8'b1111101: c <= 9'b110010110;
				8'b101001: c <= 9'b111001000;
				8'b1010010: c <= 9'b10011010;
				8'b1011000: c <= 9'b10;
				8'b101110: c <= 9'b110001111;
				8'b1000001: c <= 9'b110100;
				default: c <= 9'b0;
			endcase
			9'b110110110 : case(di)
				8'b1000011: c <= 9'b10000010;
				8'b101000: c <= 9'b110000000;
				8'b111010: c <= 9'b100111110;
				8'b110110: c <= 9'b10011011;
				8'b1100100: c <= 9'b1111011;
				8'b1000000: c <= 9'b10001001;
				8'b1110110: c <= 9'b111111111;
				8'b100101: c <= 9'b101110100;
				8'b101111: c <= 9'b110000001;
				8'b100110: c <= 9'b100100110;
				8'b1100011: c <= 9'b10100110;
				8'b1001000: c <= 9'b101000110;
				8'b111000: c <= 9'b11110001;
				8'b110001: c <= 9'b1100010;
				8'b1010111: c <= 9'b101110001;
				8'b1001110: c <= 9'b111011110;
				8'b1101010: c <= 9'b101110011;
				8'b1001001: c <= 9'b110100100;
				8'b1100000: c <= 9'b101001100;
				8'b110111: c <= 9'b101110001;
				8'b1011101: c <= 9'b101000011;
				8'b1011011: c <= 9'b110000111;
				8'b111001: c <= 9'b10101111;
				8'b1001010: c <= 9'b111111001;
				8'b110011: c <= 9'b10011101;
				8'b1101100: c <= 9'b100010101;
				8'b1110111: c <= 9'b111010110;
				8'b101011: c <= 9'b11000110;
				8'b1101011: c <= 9'b10111010;
				8'b111100: c <= 9'b111011111;
				8'b1000111: c <= 9'b111101111;
				8'b1011111: c <= 9'b110101100;
				8'b1110100: c <= 9'b100101;
				8'b101101: c <= 9'b111010000;
				8'b1010011: c <= 9'b10010;
				8'b1100001: c <= 9'b111;
				8'b110101: c <= 9'b101110100;
				8'b1000100: c <= 9'b111110000;
				8'b1010001: c <= 9'b1100001;
				8'b1010100: c <= 9'b10100011;
				8'b1100110: c <= 9'b111001001;
				8'b101010: c <= 9'b110100110;
				8'b1011110: c <= 9'b10;
				8'b1100111: c <= 9'b110001100;
				8'b1011010: c <= 9'b1010101;
				8'b1000010: c <= 9'b10100010;
				8'b111101: c <= 9'b10101011;
				8'b110000: c <= 9'b111001010;
				8'b111110: c <= 9'b101011101;
				8'b1100010: c <= 9'b110001011;
				8'b1110000: c <= 9'b110110101;
				8'b1101001: c <= 9'b100101111;
				8'b1110011: c <= 9'b11000001;
				8'b1001100: c <= 9'b110011011;
				8'b100001: c <= 9'b110110101;
				8'b1000110: c <= 9'b110001111;
				8'b1110010: c <= 9'b100000001;
				8'b1010000: c <= 9'b11011001;
				8'b1111010: c <= 9'b100001101;
				8'b1010101: c <= 9'b110101110;
				8'b111011: c <= 9'b100010;
				8'b1001101: c <= 9'b11010111;
				8'b111111: c <= 9'b111111011;
				8'b1101110: c <= 9'b110101010;
				8'b1111011: c <= 9'b100000111;
				8'b1001011: c <= 9'b10111100;
				8'b1101111: c <= 9'b1100011;
				8'b1101000: c <= 9'b1011110;
				8'b101100: c <= 9'b1000010;
				8'b100100: c <= 9'b10011010;
				8'b1111000: c <= 9'b101011101;
				8'b1000101: c <= 9'b1000100;
				8'b1011001: c <= 9'b11110111;
				8'b110100: c <= 9'b1001111;
				8'b1111001: c <= 9'b10101010;
				8'b1110001: c <= 9'b101100001;
				8'b1001111: c <= 9'b10001100;
				8'b1100101: c <= 9'b110010101;
				8'b1111110: c <= 9'b111100010;
				8'b1111100: c <= 9'b101000100;
				8'b1010110: c <= 9'b101011011;
				8'b110010: c <= 9'b100100101;
				8'b1101101: c <= 9'b100001;
				8'b100011: c <= 9'b1110;
				8'b1110101: c <= 9'b100110100;
				8'b1111101: c <= 9'b111110001;
				8'b101001: c <= 9'b11110;
				8'b1010010: c <= 9'b111001111;
				8'b1011000: c <= 9'b111111000;
				8'b101110: c <= 9'b100011;
				8'b1000001: c <= 9'b11011101;
				default: c <= 9'b0;
			endcase
			9'b101000010 : case(di)
				8'b1000011: c <= 9'b110000110;
				8'b101000: c <= 9'b111101;
				8'b111010: c <= 9'b111001000;
				8'b110110: c <= 9'b100111101;
				8'b1100100: c <= 9'b100101111;
				8'b1000000: c <= 9'b101100011;
				8'b1110110: c <= 9'b110111001;
				8'b100101: c <= 9'b100010100;
				8'b101111: c <= 9'b110111000;
				8'b100110: c <= 9'b11101101;
				8'b1100011: c <= 9'b10001010;
				8'b1001000: c <= 9'b101110;
				8'b111000: c <= 9'b100111011;
				8'b110001: c <= 9'b101010101;
				8'b1010111: c <= 9'b11000001;
				8'b1001110: c <= 9'b111010100;
				8'b1101010: c <= 9'b10011;
				8'b1001001: c <= 9'b110111011;
				8'b1100000: c <= 9'b10001110;
				8'b110111: c <= 9'b100111101;
				8'b1011101: c <= 9'b101100110;
				8'b1011011: c <= 9'b11100;
				8'b111001: c <= 9'b110000011;
				8'b1001010: c <= 9'b101010011;
				8'b110011: c <= 9'b101101100;
				8'b1101100: c <= 9'b1110000;
				8'b1110111: c <= 9'b100110100;
				8'b101011: c <= 9'b110011010;
				8'b1101011: c <= 9'b10;
				8'b111100: c <= 9'b10110100;
				8'b1000111: c <= 9'b11100001;
				8'b1011111: c <= 9'b1111110;
				8'b1110100: c <= 9'b101001010;
				8'b101101: c <= 9'b1000111;
				8'b1010011: c <= 9'b101010110;
				8'b1100001: c <= 9'b1010101;
				8'b110101: c <= 9'b101011011;
				8'b1000100: c <= 9'b101110;
				8'b1010001: c <= 9'b100110101;
				8'b1010100: c <= 9'b10101000;
				8'b1100110: c <= 9'b11111001;
				8'b101010: c <= 9'b10001100;
				8'b1011110: c <= 9'b10011001;
				8'b1100111: c <= 9'b110100;
				8'b1011010: c <= 9'b110101001;
				8'b1000010: c <= 9'b101011010;
				8'b111101: c <= 9'b100111101;
				8'b110000: c <= 9'b100101001;
				8'b111110: c <= 9'b10100011;
				8'b1100010: c <= 9'b100100011;
				8'b1110000: c <= 9'b1011;
				8'b1101001: c <= 9'b10101101;
				8'b1110011: c <= 9'b101011101;
				8'b1001100: c <= 9'b100101011;
				8'b100001: c <= 9'b100111011;
				8'b1000110: c <= 9'b101110000;
				8'b1110010: c <= 9'b1000100;
				8'b1010000: c <= 9'b11001;
				8'b1111010: c <= 9'b111100101;
				8'b1010101: c <= 9'b1111010;
				8'b111011: c <= 9'b101110010;
				8'b1001101: c <= 9'b110010010;
				8'b111111: c <= 9'b11011001;
				8'b1101110: c <= 9'b11001101;
				8'b1111011: c <= 9'b111101101;
				8'b1001011: c <= 9'b110000010;
				8'b1101111: c <= 9'b110001111;
				8'b1101000: c <= 9'b101111000;
				8'b101100: c <= 9'b10111101;
				8'b100100: c <= 9'b11001;
				8'b1111000: c <= 9'b101101010;
				8'b1000101: c <= 9'b1101;
				8'b1011001: c <= 9'b101001110;
				8'b110100: c <= 9'b100010010;
				8'b1111001: c <= 9'b10100101;
				8'b1110001: c <= 9'b10111000;
				8'b1001111: c <= 9'b110011111;
				8'b1100101: c <= 9'b111001001;
				8'b1111110: c <= 9'b100010111;
				8'b1111100: c <= 9'b100001001;
				8'b1010110: c <= 9'b11110000;
				8'b110010: c <= 9'b110011001;
				8'b1101101: c <= 9'b101;
				8'b100011: c <= 9'b111001001;
				8'b1110101: c <= 9'b11100011;
				8'b1111101: c <= 9'b10010101;
				8'b101001: c <= 9'b101110100;
				8'b1010010: c <= 9'b1111000;
				8'b1011000: c <= 9'b101110101;
				8'b101110: c <= 9'b110111110;
				8'b1000001: c <= 9'b101000100;
				default: c <= 9'b0;
			endcase
			9'b10001110 : case(di)
				8'b1000011: c <= 9'b101000010;
				8'b101000: c <= 9'b10101000;
				8'b111010: c <= 9'b11111001;
				8'b110110: c <= 9'b10110;
				8'b1100100: c <= 9'b11111010;
				8'b1000000: c <= 9'b100111100;
				8'b1110110: c <= 9'b1011010;
				8'b100101: c <= 9'b1001001;
				8'b101111: c <= 9'b10011100;
				8'b100110: c <= 9'b101110110;
				8'b1100011: c <= 9'b100100011;
				8'b1001000: c <= 9'b111000110;
				8'b111000: c <= 9'b1110001;
				8'b110001: c <= 9'b11101001;
				8'b1010111: c <= 9'b110101110;
				8'b1001110: c <= 9'b100010101;
				8'b1101010: c <= 9'b1000011;
				8'b1001001: c <= 9'b100001110;
				8'b1100000: c <= 9'b11100;
				8'b110111: c <= 9'b1111010;
				8'b1011101: c <= 9'b100001001;
				8'b1011011: c <= 9'b100000011;
				8'b111001: c <= 9'b1100011;
				8'b1001010: c <= 9'b101010110;
				8'b110011: c <= 9'b10110101;
				8'b1101100: c <= 9'b110011;
				8'b1110111: c <= 9'b101111000;
				8'b101011: c <= 9'b10010001;
				8'b1101011: c <= 9'b1010101;
				8'b111100: c <= 9'b100111001;
				8'b1000111: c <= 9'b10111101;
				8'b1011111: c <= 9'b100000110;
				8'b1110100: c <= 9'b110101111;
				8'b101101: c <= 9'b10100100;
				8'b1010011: c <= 9'b11001001;
				8'b1100001: c <= 9'b111000011;
				8'b110101: c <= 9'b100110;
				8'b1000100: c <= 9'b10;
				8'b1010001: c <= 9'b11100101;
				8'b1010100: c <= 9'b11101;
				8'b1100110: c <= 9'b10111001;
				8'b101010: c <= 9'b11001101;
				8'b1011110: c <= 9'b100110111;
				8'b1100111: c <= 9'b11110111;
				8'b1011010: c <= 9'b11100111;
				8'b1000010: c <= 9'b11001101;
				8'b111101: c <= 9'b110100001;
				8'b110000: c <= 9'b11000011;
				8'b111110: c <= 9'b1000011;
				8'b1100010: c <= 9'b110010010;
				8'b1110000: c <= 9'b110100101;
				8'b1101001: c <= 9'b100111100;
				8'b1110011: c <= 9'b101110001;
				8'b1001100: c <= 9'b110111100;
				8'b100001: c <= 9'b11001001;
				8'b1000110: c <= 9'b10100010;
				8'b1110010: c <= 9'b110001100;
				8'b1010000: c <= 9'b1100001;
				8'b1111010: c <= 9'b11110101;
				8'b1010101: c <= 9'b110000000;
				8'b111011: c <= 9'b10000010;
				8'b1001101: c <= 9'b100010010;
				8'b111111: c <= 9'b1110101;
				8'b1101110: c <= 9'b111000;
				8'b1111011: c <= 9'b100011001;
				8'b1001011: c <= 9'b11011101;
				8'b1101111: c <= 9'b1001000;
				8'b1101000: c <= 9'b111000101;
				8'b101100: c <= 9'b110000111;
				8'b100100: c <= 9'b110101011;
				8'b1111000: c <= 9'b10101;
				8'b1000101: c <= 9'b100001111;
				8'b1011001: c <= 9'b100011000;
				8'b110100: c <= 9'b1010111;
				8'b1111001: c <= 9'b11;
				8'b1110001: c <= 9'b110011001;
				8'b1001111: c <= 9'b101000101;
				8'b1100101: c <= 9'b1100101;
				8'b1111110: c <= 9'b101001;
				8'b1111100: c <= 9'b111100001;
				8'b1010110: c <= 9'b100000001;
				8'b110010: c <= 9'b11101000;
				8'b1101101: c <= 9'b111000000;
				8'b100011: c <= 9'b111000011;
				8'b1110101: c <= 9'b110010010;
				8'b1111101: c <= 9'b111111;
				8'b101001: c <= 9'b1010010;
				8'b1010010: c <= 9'b10011111;
				8'b1011000: c <= 9'b101101100;
				8'b101110: c <= 9'b10010100;
				8'b1000001: c <= 9'b10101010;
				default: c <= 9'b0;
			endcase
			9'b11111010 : case(di)
				8'b1000011: c <= 9'b1011000;
				8'b101000: c <= 9'b100111101;
				8'b111010: c <= 9'b1101111;
				8'b110110: c <= 9'b100101001;
				8'b1100100: c <= 9'b111001010;
				8'b1000000: c <= 9'b110010;
				8'b1110110: c <= 9'b101000100;
				8'b100101: c <= 9'b111000110;
				8'b101111: c <= 9'b101000111;
				8'b100110: c <= 9'b1011;
				8'b1100011: c <= 9'b111011110;
				8'b1001000: c <= 9'b111001010;
				8'b111000: c <= 9'b11110100;
				8'b110001: c <= 9'b100010100;
				8'b1010111: c <= 9'b111101001;
				8'b1001110: c <= 9'b101011111;
				8'b1101010: c <= 9'b111110110;
				8'b1001001: c <= 9'b100001010;
				8'b1100000: c <= 9'b111010000;
				8'b110111: c <= 9'b11010;
				8'b1011101: c <= 9'b1101111;
				8'b1011011: c <= 9'b11010001;
				8'b111001: c <= 9'b101110000;
				8'b1001010: c <= 9'b100101001;
				8'b110011: c <= 9'b111110101;
				8'b1101100: c <= 9'b101011;
				8'b1110111: c <= 9'b11111010;
				8'b101011: c <= 9'b100000110;
				8'b1101011: c <= 9'b101110001;
				8'b111100: c <= 9'b10000011;
				8'b1000111: c <= 9'b10100;
				8'b1011111: c <= 9'b111100111;
				8'b1110100: c <= 9'b10010110;
				8'b101101: c <= 9'b101110000;
				8'b1010011: c <= 9'b10001010;
				8'b1100001: c <= 9'b1000110;
				8'b110101: c <= 9'b1011001;
				8'b1000100: c <= 9'b1011111;
				8'b1010001: c <= 9'b1010001;
				8'b1010100: c <= 9'b11100;
				8'b1100110: c <= 9'b111111101;
				8'b101010: c <= 9'b111111000;
				8'b1011110: c <= 9'b11110010;
				8'b1100111: c <= 9'b10101000;
				8'b1011010: c <= 9'b100010001;
				8'b1000010: c <= 9'b101000011;
				8'b111101: c <= 9'b100110;
				8'b110000: c <= 9'b11001001;
				8'b111110: c <= 9'b10001000;
				8'b1100010: c <= 9'b100000000;
				8'b1110000: c <= 9'b11001111;
				8'b1101001: c <= 9'b1001110;
				8'b1110011: c <= 9'b10101;
				8'b1001100: c <= 9'b11111011;
				8'b100001: c <= 9'b10101;
				8'b1000110: c <= 9'b101000011;
				8'b1110010: c <= 9'b100001111;
				8'b1010000: c <= 9'b11100110;
				8'b1111010: c <= 9'b111;
				8'b1010101: c <= 9'b110000011;
				8'b111011: c <= 9'b1000001;
				8'b1001101: c <= 9'b110010101;
				8'b111111: c <= 9'b111110110;
				8'b1101110: c <= 9'b10111000;
				8'b1111011: c <= 9'b10111011;
				8'b1001011: c <= 9'b1111000;
				8'b1101111: c <= 9'b10000;
				8'b1101000: c <= 9'b110111;
				8'b101100: c <= 9'b1011000;
				8'b100100: c <= 9'b101101100;
				8'b1111000: c <= 9'b11111010;
				8'b1000101: c <= 9'b10011101;
				8'b1011001: c <= 9'b111000010;
				8'b110100: c <= 9'b100011000;
				8'b1111001: c <= 9'b101010001;
				8'b1110001: c <= 9'b100101110;
				8'b1001111: c <= 9'b110111;
				8'b1100101: c <= 9'b1100001;
				8'b1111110: c <= 9'b1010001;
				8'b1111100: c <= 9'b11100;
				8'b1010110: c <= 9'b11001011;
				8'b110010: c <= 9'b11001001;
				8'b1101101: c <= 9'b101100010;
				8'b100011: c <= 9'b100101110;
				8'b1110101: c <= 9'b10001110;
				8'b1111101: c <= 9'b10000010;
				8'b101001: c <= 9'b110001010;
				8'b1010010: c <= 9'b100110111;
				8'b1011000: c <= 9'b1101001;
				8'b101110: c <= 9'b111001100;
				8'b1000001: c <= 9'b111010111;
				default: c <= 9'b0;
			endcase
			9'b110100001 : case(di)
				8'b1000011: c <= 9'b111001100;
				8'b101000: c <= 9'b110001110;
				8'b111010: c <= 9'b101110010;
				8'b110110: c <= 9'b100010001;
				8'b1100100: c <= 9'b100010100;
				8'b1000000: c <= 9'b11100010;
				8'b1110110: c <= 9'b110100100;
				8'b100101: c <= 9'b101001110;
				8'b101111: c <= 9'b10010110;
				8'b100110: c <= 9'b11001010;
				8'b1100011: c <= 9'b100100101;
				8'b1001000: c <= 9'b11111011;
				8'b111000: c <= 9'b100011001;
				8'b110001: c <= 9'b1000101;
				8'b1010111: c <= 9'b10111000;
				8'b1001110: c <= 9'b11101100;
				8'b1101010: c <= 9'b101010001;
				8'b1001001: c <= 9'b10010111;
				8'b1100000: c <= 9'b101110100;
				8'b110111: c <= 9'b110010;
				8'b1011101: c <= 9'b100011;
				8'b1011011: c <= 9'b111011111;
				8'b111001: c <= 9'b101000010;
				8'b1001010: c <= 9'b1001100;
				8'b110011: c <= 9'b101001111;
				8'b1101100: c <= 9'b110110010;
				8'b1110111: c <= 9'b1011111;
				8'b101011: c <= 9'b111001011;
				8'b1101011: c <= 9'b111010111;
				8'b111100: c <= 9'b11100101;
				8'b1000111: c <= 9'b10110100;
				8'b1011111: c <= 9'b1111101;
				8'b1110100: c <= 9'b10101100;
				8'b101101: c <= 9'b101110001;
				8'b1010011: c <= 9'b1111;
				8'b1100001: c <= 9'b100001001;
				8'b110101: c <= 9'b11110;
				8'b1000100: c <= 9'b101110111;
				8'b1010001: c <= 9'b1001111;
				8'b1010100: c <= 9'b100100111;
				8'b1100110: c <= 9'b100001111;
				8'b101010: c <= 9'b11010101;
				8'b1011110: c <= 9'b101100101;
				8'b1100111: c <= 9'b10100111;
				8'b1011010: c <= 9'b1111010;
				8'b1000010: c <= 9'b10110;
				8'b111101: c <= 9'b11111000;
				8'b110000: c <= 9'b101011101;
				8'b111110: c <= 9'b101100111;
				8'b1100010: c <= 9'b101100000;
				8'b1110000: c <= 9'b111001;
				8'b1101001: c <= 9'b10000101;
				8'b1110011: c <= 9'b111001011;
				8'b1001100: c <= 9'b1010010;
				8'b100001: c <= 9'b111100001;
				8'b1000110: c <= 9'b111111010;
				8'b1110010: c <= 9'b1101001;
				8'b1010000: c <= 9'b111000011;
				8'b1111010: c <= 9'b111001001;
				8'b1010101: c <= 9'b10100111;
				8'b111011: c <= 9'b1001000;
				8'b1001101: c <= 9'b111011001;
				8'b111111: c <= 9'b11101;
				8'b1101110: c <= 9'b110000101;
				8'b1111011: c <= 9'b10111010;
				8'b1001011: c <= 9'b110010111;
				8'b1101111: c <= 9'b111011101;
				8'b1101000: c <= 9'b110110;
				8'b101100: c <= 9'b11001110;
				8'b100100: c <= 9'b111011100;
				8'b1111000: c <= 9'b1110100;
				8'b1000101: c <= 9'b1001110;
				8'b1011001: c <= 9'b101000110;
				8'b110100: c <= 9'b11001010;
				8'b1111001: c <= 9'b11100010;
				8'b1110001: c <= 9'b11100101;
				8'b1001111: c <= 9'b111101;
				8'b1100101: c <= 9'b1101;
				8'b1111110: c <= 9'b111111111;
				8'b1111100: c <= 9'b11100101;
				8'b1010110: c <= 9'b101110110;
				8'b110010: c <= 9'b11101000;
				8'b1101101: c <= 9'b1011111;
				8'b100011: c <= 9'b10010111;
				8'b1110101: c <= 9'b101000001;
				8'b1111101: c <= 9'b101111000;
				8'b101001: c <= 9'b1001100;
				8'b1010010: c <= 9'b100110011;
				8'b1011000: c <= 9'b110001010;
				8'b101110: c <= 9'b111010;
				8'b1000001: c <= 9'b110110010;
				default: c <= 9'b0;
			endcase
			9'b100100000 : case(di)
				8'b1000011: c <= 9'b1000001;
				8'b101000: c <= 9'b111101100;
				8'b111010: c <= 9'b100111001;
				8'b110110: c <= 9'b1001000;
				8'b1100100: c <= 9'b101001011;
				8'b1000000: c <= 9'b110001111;
				8'b1110110: c <= 9'b111100110;
				8'b100101: c <= 9'b110011100;
				8'b101111: c <= 9'b1001010;
				8'b100110: c <= 9'b10001001;
				8'b1100011: c <= 9'b110111001;
				8'b1001000: c <= 9'b100100110;
				8'b111000: c <= 9'b100011101;
				8'b110001: c <= 9'b10100000;
				8'b1010111: c <= 9'b111011;
				8'b1001110: c <= 9'b1000101;
				8'b1101010: c <= 9'b1001000;
				8'b1001001: c <= 9'b1010011;
				8'b1100000: c <= 9'b110011000;
				8'b110111: c <= 9'b111001110;
				8'b1011101: c <= 9'b10111101;
				8'b1011011: c <= 9'b10101;
				8'b111001: c <= 9'b111111000;
				8'b1001010: c <= 9'b10111001;
				8'b110011: c <= 9'b111101000;
				8'b1101100: c <= 9'b10;
				8'b1110111: c <= 9'b11001100;
				8'b101011: c <= 9'b1100;
				8'b1101011: c <= 9'b101101111;
				8'b111100: c <= 9'b11000011;
				8'b1000111: c <= 9'b101110100;
				8'b1011111: c <= 9'b10010111;
				8'b1110100: c <= 9'b11001;
				8'b101101: c <= 9'b11110001;
				8'b1010011: c <= 9'b11100110;
				8'b1100001: c <= 9'b10011000;
				8'b110101: c <= 9'b111100101;
				8'b1000100: c <= 9'b111101010;
				8'b1010001: c <= 9'b101011111;
				8'b1010100: c <= 9'b101100111;
				8'b1100110: c <= 9'b11001100;
				8'b101010: c <= 9'b1111100;
				8'b1011110: c <= 9'b11000111;
				8'b1100111: c <= 9'b11010101;
				8'b1011010: c <= 9'b11010010;
				8'b1000010: c <= 9'b100001110;
				8'b111101: c <= 9'b101110100;
				8'b110000: c <= 9'b101001000;
				8'b111110: c <= 9'b100101011;
				8'b1100010: c <= 9'b100011010;
				8'b1110000: c <= 9'b100001;
				8'b1101001: c <= 9'b11011000;
				8'b1110011: c <= 9'b110000111;
				8'b1001100: c <= 9'b11000110;
				8'b100001: c <= 9'b11011001;
				8'b1000110: c <= 9'b11111100;
				8'b1110010: c <= 9'b110101111;
				8'b1010000: c <= 9'b100011011;
				8'b1111010: c <= 9'b11100010;
				8'b1010101: c <= 9'b101111111;
				8'b111011: c <= 9'b110101011;
				8'b1001101: c <= 9'b11110000;
				8'b111111: c <= 9'b101100000;
				8'b1101110: c <= 9'b11111011;
				8'b1111011: c <= 9'b11110010;
				8'b1001011: c <= 9'b101011;
				8'b1101111: c <= 9'b110010101;
				8'b1101000: c <= 9'b1010010;
				8'b101100: c <= 9'b111101;
				8'b100100: c <= 9'b10111110;
				8'b1111000: c <= 9'b11101101;
				8'b1000101: c <= 9'b1111011;
				8'b1011001: c <= 9'b101001011;
				8'b110100: c <= 9'b100100;
				8'b1111001: c <= 9'b100001110;
				8'b1110001: c <= 9'b111011101;
				8'b1001111: c <= 9'b11011010;
				8'b1100101: c <= 9'b100001100;
				8'b1111110: c <= 9'b10110101;
				8'b1111100: c <= 9'b11110111;
				8'b1010110: c <= 9'b1111101;
				8'b110010: c <= 9'b110011010;
				8'b1101101: c <= 9'b100101101;
				8'b100011: c <= 9'b11101011;
				8'b1110101: c <= 9'b10111000;
				8'b1111101: c <= 9'b101000010;
				8'b101001: c <= 9'b10001110;
				8'b1010010: c <= 9'b1110011;
				8'b1011000: c <= 9'b110000;
				8'b101110: c <= 9'b1100100;
				8'b1000001: c <= 9'b1100101;
				default: c <= 9'b0;
			endcase
			9'b111001111 : case(di)
				8'b1000011: c <= 9'b101110101;
				8'b101000: c <= 9'b11101000;
				8'b111010: c <= 9'b11010001;
				8'b110110: c <= 9'b1000111;
				8'b1100100: c <= 9'b101100111;
				8'b1000000: c <= 9'b110100001;
				8'b1110110: c <= 9'b101111000;
				8'b100101: c <= 9'b1101101;
				8'b101111: c <= 9'b110110;
				8'b100110: c <= 9'b11011;
				8'b1100011: c <= 9'b110001000;
				8'b1001000: c <= 9'b100110100;
				8'b111000: c <= 9'b110110011;
				8'b110001: c <= 9'b10101;
				8'b1010111: c <= 9'b111000011;
				8'b1001110: c <= 9'b101101000;
				8'b1101010: c <= 9'b110111000;
				8'b1001001: c <= 9'b111010000;
				8'b1100000: c <= 9'b10111101;
				8'b110111: c <= 9'b111100000;
				8'b1011101: c <= 9'b110111001;
				8'b1011011: c <= 9'b1000001;
				8'b111001: c <= 9'b110011000;
				8'b1001010: c <= 9'b110111000;
				8'b110011: c <= 9'b111011010;
				8'b1101100: c <= 9'b101101110;
				8'b1110111: c <= 9'b110011011;
				8'b101011: c <= 9'b101101111;
				8'b1101011: c <= 9'b11011100;
				8'b111100: c <= 9'b101001010;
				8'b1000111: c <= 9'b1011000;
				8'b1011111: c <= 9'b110011;
				8'b1110100: c <= 9'b11111011;
				8'b101101: c <= 9'b11101111;
				8'b1010011: c <= 9'b1001100;
				8'b1100001: c <= 9'b100001110;
				8'b110101: c <= 9'b1000111;
				8'b1000100: c <= 9'b101001000;
				8'b1010001: c <= 9'b1100;
				8'b1010100: c <= 9'b111101;
				8'b1100110: c <= 9'b10100011;
				8'b101010: c <= 9'b100011111;
				8'b1011110: c <= 9'b11100010;
				8'b1100111: c <= 9'b110001111;
				8'b1011010: c <= 9'b11010011;
				8'b1000010: c <= 9'b100000100;
				8'b111101: c <= 9'b100011;
				8'b110000: c <= 9'b11100101;
				8'b111110: c <= 9'b101011011;
				8'b1100010: c <= 9'b1011;
				8'b1110000: c <= 9'b1110101;
				8'b1101001: c <= 9'b10000110;
				8'b1110011: c <= 9'b100111111;
				8'b1001100: c <= 9'b10011111;
				8'b100001: c <= 9'b111100000;
				8'b1000110: c <= 9'b110111010;
				8'b1110010: c <= 9'b11110;
				8'b1010000: c <= 9'b101101000;
				8'b1111010: c <= 9'b100101100;
				8'b1010101: c <= 9'b10101101;
				8'b111011: c <= 9'b100001001;
				8'b1001101: c <= 9'b10011010;
				8'b111111: c <= 9'b110111111;
				8'b1101110: c <= 9'b11001100;
				8'b1111011: c <= 9'b11100;
				8'b1001011: c <= 9'b10100101;
				8'b1101111: c <= 9'b111011111;
				8'b1101000: c <= 9'b101010011;
				8'b101100: c <= 9'b110100010;
				8'b100100: c <= 9'b100101011;
				8'b1111000: c <= 9'b101111110;
				8'b1000101: c <= 9'b10001000;
				8'b1011001: c <= 9'b100001110;
				8'b110100: c <= 9'b11011000;
				8'b1111001: c <= 9'b1101;
				8'b1110001: c <= 9'b11011010;
				8'b1001111: c <= 9'b11011001;
				8'b1100101: c <= 9'b111100110;
				8'b1111110: c <= 9'b100110011;
				8'b1111100: c <= 9'b100001110;
				8'b1010110: c <= 9'b1100011;
				8'b110010: c <= 9'b100101001;
				8'b1101101: c <= 9'b10111000;
				8'b100011: c <= 9'b111000110;
				8'b1110101: c <= 9'b1011010;
				8'b1111101: c <= 9'b111100111;
				8'b101001: c <= 9'b101110011;
				8'b1010010: c <= 9'b10100101;
				8'b1011000: c <= 9'b1110001;
				8'b101110: c <= 9'b11101101;
				8'b1000001: c <= 9'b10110010;
				default: c <= 9'b0;
			endcase
			9'b110101100 : case(di)
				8'b1000011: c <= 9'b101110100;
				8'b101000: c <= 9'b100010000;
				8'b111010: c <= 9'b100011100;
				8'b110110: c <= 9'b110111011;
				8'b1100100: c <= 9'b10011000;
				8'b1000000: c <= 9'b100001010;
				8'b1110110: c <= 9'b1010101;
				8'b100101: c <= 9'b10011101;
				8'b101111: c <= 9'b11110100;
				8'b100110: c <= 9'b111011;
				8'b1100011: c <= 9'b1010000;
				8'b1001000: c <= 9'b101010101;
				8'b111000: c <= 9'b110011011;
				8'b110001: c <= 9'b11101;
				8'b1010111: c <= 9'b111010100;
				8'b1001110: c <= 9'b10011101;
				8'b1101010: c <= 9'b100100011;
				8'b1001001: c <= 9'b110100010;
				8'b1100000: c <= 9'b1001011;
				8'b110111: c <= 9'b1001101;
				8'b1011101: c <= 9'b111000110;
				8'b1011011: c <= 9'b10;
				8'b111001: c <= 9'b101101011;
				8'b1001010: c <= 9'b111001100;
				8'b110011: c <= 9'b111011;
				8'b1101100: c <= 9'b110000;
				8'b1110111: c <= 9'b101100010;
				8'b101011: c <= 9'b11111;
				8'b1101011: c <= 9'b10101;
				8'b111100: c <= 9'b11100;
				8'b1000111: c <= 9'b100100;
				8'b1011111: c <= 9'b100000110;
				8'b1110100: c <= 9'b10101111;
				8'b101101: c <= 9'b100111010;
				8'b1010011: c <= 9'b100100;
				8'b1100001: c <= 9'b1100000;
				8'b110101: c <= 9'b1011010;
				8'b1000100: c <= 9'b11010111;
				8'b1010001: c <= 9'b110110010;
				8'b1010100: c <= 9'b110110111;
				8'b1100110: c <= 9'b111111001;
				8'b101010: c <= 9'b100000001;
				8'b1011110: c <= 9'b110100111;
				8'b1100111: c <= 9'b11000111;
				8'b1011010: c <= 9'b110010;
				8'b1000010: c <= 9'b110100110;
				8'b111101: c <= 9'b101100001;
				8'b110000: c <= 9'b101001100;
				8'b111110: c <= 9'b10011001;
				8'b1100010: c <= 9'b110111000;
				8'b1110000: c <= 9'b10110101;
				8'b1101001: c <= 9'b10100110;
				8'b1110011: c <= 9'b100111011;
				8'b1001100: c <= 9'b111011100;
				8'b100001: c <= 9'b110100110;
				8'b1000110: c <= 9'b110111011;
				8'b1110010: c <= 9'b110111110;
				8'b1010000: c <= 9'b111000110;
				8'b1111010: c <= 9'b100011010;
				8'b1010101: c <= 9'b100100;
				8'b111011: c <= 9'b100100011;
				8'b1001101: c <= 9'b110001000;
				8'b111111: c <= 9'b100010111;
				8'b1101110: c <= 9'b100010100;
				8'b1111011: c <= 9'b100011010;
				8'b1001011: c <= 9'b101001100;
				8'b1101111: c <= 9'b101111010;
				8'b1101000: c <= 9'b100110110;
				8'b101100: c <= 9'b11100010;
				8'b100100: c <= 9'b110100000;
				8'b1111000: c <= 9'b1000111;
				8'b1000101: c <= 9'b1011001;
				8'b1011001: c <= 9'b101110011;
				8'b110100: c <= 9'b101110011;
				8'b1111001: c <= 9'b100010;
				8'b1110001: c <= 9'b100000000;
				8'b1001111: c <= 9'b101101011;
				8'b1100101: c <= 9'b110000010;
				8'b1111110: c <= 9'b110100011;
				8'b1111100: c <= 9'b1000110;
				8'b1010110: c <= 9'b111010;
				8'b110010: c <= 9'b101010011;
				8'b1101101: c <= 9'b10101100;
				8'b100011: c <= 9'b100010100;
				8'b1110101: c <= 9'b100001010;
				8'b1111101: c <= 9'b101011;
				8'b101001: c <= 9'b110010010;
				8'b1010010: c <= 9'b1100100;
				8'b1011000: c <= 9'b10000010;
				8'b101110: c <= 9'b11111001;
				8'b1000001: c <= 9'b11100001;
				default: c <= 9'b0;
			endcase
			9'b10110101 : case(di)
				8'b1000011: c <= 9'b11101000;
				8'b101000: c <= 9'b1101;
				8'b111010: c <= 9'b110011010;
				8'b110110: c <= 9'b100100010;
				8'b1100100: c <= 9'b11001111;
				8'b1000000: c <= 9'b101000110;
				8'b1110110: c <= 9'b10110001;
				8'b100101: c <= 9'b1101101;
				8'b101111: c <= 9'b110101011;
				8'b100110: c <= 9'b1100011;
				8'b1100011: c <= 9'b11110110;
				8'b1001000: c <= 9'b101110110;
				8'b111000: c <= 9'b101001;
				8'b110001: c <= 9'b100000000;
				8'b1010111: c <= 9'b11001110;
				8'b1001110: c <= 9'b101111010;
				8'b1101010: c <= 9'b111101100;
				8'b1001001: c <= 9'b111100011;
				8'b1100000: c <= 9'b110001;
				8'b110111: c <= 9'b111101111;
				8'b1011101: c <= 9'b1101000;
				8'b1011011: c <= 9'b110101;
				8'b111001: c <= 9'b11011;
				8'b1001010: c <= 9'b10000;
				8'b110011: c <= 9'b1011001;
				8'b1101100: c <= 9'b1111000;
				8'b1110111: c <= 9'b111111010;
				8'b101011: c <= 9'b100110110;
				8'b1101011: c <= 9'b11111001;
				8'b111100: c <= 9'b101001111;
				8'b1000111: c <= 9'b11111110;
				8'b1011111: c <= 9'b1000;
				8'b1110100: c <= 9'b101111111;
				8'b101101: c <= 9'b1001001;
				8'b1010011: c <= 9'b101010001;
				8'b1100001: c <= 9'b100101111;
				8'b110101: c <= 9'b10110001;
				8'b1000100: c <= 9'b100000110;
				8'b1010001: c <= 9'b1111100;
				8'b1010100: c <= 9'b10100010;
				8'b1100110: c <= 9'b11010000;
				8'b101010: c <= 9'b10;
				8'b1011110: c <= 9'b111101001;
				8'b1100111: c <= 9'b100110011;
				8'b1011010: c <= 9'b11110;
				8'b1000010: c <= 9'b1001001;
				8'b111101: c <= 9'b110101100;
				8'b110000: c <= 9'b10010000;
				8'b111110: c <= 9'b1001001;
				8'b1100010: c <= 9'b11011;
				8'b1110000: c <= 9'b1101111;
				8'b1101001: c <= 9'b11001111;
				8'b1110011: c <= 9'b110;
				8'b1001100: c <= 9'b11010011;
				8'b100001: c <= 9'b110010011;
				8'b1000110: c <= 9'b10101010;
				8'b1110010: c <= 9'b110011011;
				8'b1010000: c <= 9'b111001010;
				8'b1111010: c <= 9'b10101110;
				8'b1010101: c <= 9'b10110101;
				8'b111011: c <= 9'b100101100;
				8'b1001101: c <= 9'b100000001;
				8'b111111: c <= 9'b100101110;
				8'b1101110: c <= 9'b111100001;
				8'b1111011: c <= 9'b101100;
				8'b1001011: c <= 9'b110110;
				8'b1101111: c <= 9'b101101011;
				8'b1101000: c <= 9'b111110001;
				8'b101100: c <= 9'b10011101;
				8'b100100: c <= 9'b101110110;
				8'b1111000: c <= 9'b10110010;
				8'b1000101: c <= 9'b100001100;
				8'b1011001: c <= 9'b10110100;
				8'b110100: c <= 9'b1001011;
				8'b1111001: c <= 9'b110011100;
				8'b1110001: c <= 9'b11100010;
				8'b1001111: c <= 9'b101011010;
				8'b1100101: c <= 9'b101010101;
				8'b1111110: c <= 9'b101100110;
				8'b1111100: c <= 9'b1110101;
				8'b1010110: c <= 9'b101101001;
				8'b110010: c <= 9'b111000000;
				8'b1101101: c <= 9'b111000000;
				8'b100011: c <= 9'b101101101;
				8'b1110101: c <= 9'b111111101;
				8'b1111101: c <= 9'b10111;
				8'b101001: c <= 9'b11000110;
				8'b1010010: c <= 9'b101000010;
				8'b1011000: c <= 9'b10010110;
				8'b101110: c <= 9'b11001010;
				8'b1000001: c <= 9'b111010010;
				default: c <= 9'b0;
			endcase
			9'b1100111 : case(di)
				8'b1000011: c <= 9'b101001111;
				8'b101000: c <= 9'b110100110;
				8'b111010: c <= 9'b111100110;
				8'b110110: c <= 9'b1111;
				8'b1100100: c <= 9'b10110111;
				8'b1000000: c <= 9'b110000110;
				8'b1110110: c <= 9'b111110001;
				8'b100101: c <= 9'b111101100;
				8'b101111: c <= 9'b10001010;
				8'b100110: c <= 9'b101011110;
				8'b1100011: c <= 9'b110010;
				8'b1001000: c <= 9'b10110;
				8'b111000: c <= 9'b10010101;
				8'b110001: c <= 9'b110110;
				8'b1010111: c <= 9'b10;
				8'b1001110: c <= 9'b111010001;
				8'b1101010: c <= 9'b111100100;
				8'b1001001: c <= 9'b1111000;
				8'b1100000: c <= 9'b100010011;
				8'b110111: c <= 9'b11011000;
				8'b1011101: c <= 9'b11001100;
				8'b1011011: c <= 9'b110111111;
				8'b111001: c <= 9'b110000111;
				8'b1001010: c <= 9'b110010001;
				8'b110011: c <= 9'b110101011;
				8'b1101100: c <= 9'b1111;
				8'b1110111: c <= 9'b10000111;
				8'b101011: c <= 9'b100010110;
				8'b1101011: c <= 9'b111010100;
				8'b111100: c <= 9'b11001011;
				8'b1000111: c <= 9'b100011111;
				8'b1011111: c <= 9'b100000110;
				8'b1110100: c <= 9'b111000010;
				8'b101101: c <= 9'b111101110;
				8'b1010011: c <= 9'b110011101;
				8'b1100001: c <= 9'b100101110;
				8'b110101: c <= 9'b1111100;
				8'b1000100: c <= 9'b110001100;
				8'b1010001: c <= 9'b11000010;
				8'b1010100: c <= 9'b101010111;
				8'b1100110: c <= 9'b11000001;
				8'b101010: c <= 9'b1110;
				8'b1011110: c <= 9'b110011001;
				8'b1100111: c <= 9'b101110111;
				8'b1011010: c <= 9'b111011110;
				8'b1000010: c <= 9'b11010101;
				8'b111101: c <= 9'b110011000;
				8'b110000: c <= 9'b100111101;
				8'b111110: c <= 9'b10010100;
				8'b1100010: c <= 9'b11111011;
				8'b1110000: c <= 9'b10100100;
				8'b1101001: c <= 9'b100110100;
				8'b1110011: c <= 9'b11110001;
				8'b1001100: c <= 9'b10110001;
				8'b100001: c <= 9'b100011;
				8'b1000110: c <= 9'b10;
				8'b1110010: c <= 9'b11001101;
				8'b1010000: c <= 9'b1100011;
				8'b1111010: c <= 9'b100111000;
				8'b1010101: c <= 9'b11011;
				8'b111011: c <= 9'b101110100;
				8'b1001101: c <= 9'b100010;
				8'b111111: c <= 9'b100101100;
				8'b1101110: c <= 9'b101011111;
				8'b1111011: c <= 9'b10110;
				8'b1001011: c <= 9'b110111010;
				8'b1101111: c <= 9'b11111010;
				8'b1101000: c <= 9'b100001100;
				8'b101100: c <= 9'b10001000;
				8'b100100: c <= 9'b100110101;
				8'b1111000: c <= 9'b100010;
				8'b1000101: c <= 9'b101101001;
				8'b1011001: c <= 9'b11001001;
				8'b110100: c <= 9'b100011111;
				8'b1111001: c <= 9'b100101000;
				8'b1110001: c <= 9'b101101111;
				8'b1001111: c <= 9'b101010011;
				8'b1100101: c <= 9'b10001111;
				8'b1111110: c <= 9'b100011100;
				8'b1111100: c <= 9'b11110011;
				8'b1010110: c <= 9'b101111001;
				8'b110010: c <= 9'b11010000;
				8'b1101101: c <= 9'b101000111;
				8'b100011: c <= 9'b111001110;
				8'b1110101: c <= 9'b11010;
				8'b1111101: c <= 9'b1000110;
				8'b101001: c <= 9'b111000000;
				8'b1010010: c <= 9'b1001100;
				8'b1011000: c <= 9'b11110010;
				8'b101110: c <= 9'b100001011;
				8'b1000001: c <= 9'b101101011;
				default: c <= 9'b0;
			endcase
			9'b110010010 : case(di)
				8'b1000011: c <= 9'b100000100;
				8'b101000: c <= 9'b11110011;
				8'b111010: c <= 9'b101010;
				8'b110110: c <= 9'b101110010;
				8'b1100100: c <= 9'b11010010;
				8'b1000000: c <= 9'b101001011;
				8'b1110110: c <= 9'b10001110;
				8'b100101: c <= 9'b1100010;
				8'b101111: c <= 9'b101110011;
				8'b100110: c <= 9'b101011010;
				8'b1100011: c <= 9'b1010111;
				8'b1001000: c <= 9'b110001001;
				8'b111000: c <= 9'b1010101;
				8'b110001: c <= 9'b111110110;
				8'b1010111: c <= 9'b1111010;
				8'b1001110: c <= 9'b11101111;
				8'b1101010: c <= 9'b1110000;
				8'b1001001: c <= 9'b1001101;
				8'b1100000: c <= 9'b110000011;
				8'b110111: c <= 9'b100011100;
				8'b1011101: c <= 9'b101001010;
				8'b1011011: c <= 9'b11110010;
				8'b111001: c <= 9'b11011000;
				8'b1001010: c <= 9'b101101111;
				8'b110011: c <= 9'b10110001;
				8'b1101100: c <= 9'b110011101;
				8'b1110111: c <= 9'b11010111;
				8'b101011: c <= 9'b100000100;
				8'b1101011: c <= 9'b111001110;
				8'b111100: c <= 9'b1000100;
				8'b1000111: c <= 9'b11010010;
				8'b1011111: c <= 9'b1100000;
				8'b1110100: c <= 9'b110110010;
				8'b101101: c <= 9'b110000101;
				8'b1010011: c <= 9'b101010001;
				8'b1100001: c <= 9'b10000001;
				8'b110101: c <= 9'b100110110;
				8'b1000100: c <= 9'b11000;
				8'b1010001: c <= 9'b101011111;
				8'b1010100: c <= 9'b110010101;
				8'b1100110: c <= 9'b100111010;
				8'b101010: c <= 9'b1101;
				8'b1011110: c <= 9'b101100101;
				8'b1100111: c <= 9'b110100001;
				8'b1011010: c <= 9'b101010100;
				8'b1000010: c <= 9'b101110111;
				8'b111101: c <= 9'b11101100;
				8'b110000: c <= 9'b101000110;
				8'b111110: c <= 9'b110101111;
				8'b1100010: c <= 9'b100101110;
				8'b1110000: c <= 9'b101001011;
				8'b1101001: c <= 9'b1000000;
				8'b1110011: c <= 9'b10111010;
				8'b1001100: c <= 9'b111011010;
				8'b100001: c <= 9'b101111110;
				8'b1000110: c <= 9'b1;
				8'b1110010: c <= 9'b100101100;
				8'b1010000: c <= 9'b1111001;
				8'b1111010: c <= 9'b1101100;
				8'b1010101: c <= 9'b11100001;
				8'b111011: c <= 9'b101010;
				8'b1001101: c <= 9'b111001110;
				8'b111111: c <= 9'b111110001;
				8'b1101110: c <= 9'b101100010;
				8'b1111011: c <= 9'b100100011;
				8'b1001011: c <= 9'b111101100;
				8'b1101111: c <= 9'b10111000;
				8'b1101000: c <= 9'b10111111;
				8'b101100: c <= 9'b111101001;
				8'b100100: c <= 9'b11010000;
				8'b1111000: c <= 9'b11101011;
				8'b1000101: c <= 9'b111100001;
				8'b1011001: c <= 9'b1101010;
				8'b110100: c <= 9'b11001000;
				8'b1111001: c <= 9'b100101000;
				8'b1110001: c <= 9'b1111010;
				8'b1001111: c <= 9'b11000000;
				8'b1100101: c <= 9'b111000101;
				8'b1111110: c <= 9'b11010001;
				8'b1111100: c <= 9'b110110100;
				8'b1010110: c <= 9'b101011101;
				8'b110010: c <= 9'b110001101;
				8'b1101101: c <= 9'b1001001;
				8'b100011: c <= 9'b10100011;
				8'b1110101: c <= 9'b111110011;
				8'b1111101: c <= 9'b1100100;
				8'b101001: c <= 9'b1111;
				8'b1010010: c <= 9'b10011101;
				8'b1011000: c <= 9'b10;
				8'b101110: c <= 9'b11111100;
				8'b1000001: c <= 9'b101010011;
				default: c <= 9'b0;
			endcase
			9'b1111101 : case(di)
				8'b1000011: c <= 9'b100011111;
				8'b101000: c <= 9'b110001100;
				8'b111010: c <= 9'b1011111;
				8'b110110: c <= 9'b110110100;
				8'b1100100: c <= 9'b11011010;
				8'b1000000: c <= 9'b101000110;
				8'b1110110: c <= 9'b111000000;
				8'b100101: c <= 9'b10001011;
				8'b101111: c <= 9'b110001110;
				8'b100110: c <= 9'b110110101;
				8'b1100011: c <= 9'b100011101;
				8'b1001000: c <= 9'b10010111;
				8'b111000: c <= 9'b10000001;
				8'b110001: c <= 9'b10100010;
				8'b1010111: c <= 9'b1011000;
				8'b1001110: c <= 9'b111110101;
				8'b1101010: c <= 9'b101010010;
				8'b1001001: c <= 9'b10001110;
				8'b1100000: c <= 9'b11;
				8'b110111: c <= 9'b111001011;
				8'b1011101: c <= 9'b1011;
				8'b1011011: c <= 9'b10100110;
				8'b111001: c <= 9'b100110110;
				8'b1001010: c <= 9'b100101000;
				8'b110011: c <= 9'b110000000;
				8'b1101100: c <= 9'b11101001;
				8'b1110111: c <= 9'b11100;
				8'b101011: c <= 9'b11000111;
				8'b1101011: c <= 9'b11100111;
				8'b111100: c <= 9'b100101110;
				8'b1000111: c <= 9'b100110101;
				8'b1011111: c <= 9'b1011011;
				8'b1110100: c <= 9'b100011101;
				8'b101101: c <= 9'b10011111;
				8'b1010011: c <= 9'b111000;
				8'b1100001: c <= 9'b11100;
				8'b110101: c <= 9'b11001000;
				8'b1000100: c <= 9'b101000101;
				8'b1010001: c <= 9'b110110101;
				8'b1010100: c <= 9'b11000000;
				8'b1100110: c <= 9'b11011010;
				8'b101010: c <= 9'b1000100;
				8'b1011110: c <= 9'b10000001;
				8'b1100111: c <= 9'b100;
				8'b1011010: c <= 9'b100111000;
				8'b1000010: c <= 9'b1011;
				8'b111101: c <= 9'b111011100;
				8'b110000: c <= 9'b101111111;
				8'b111110: c <= 9'b1100111;
				8'b1100010: c <= 9'b1111111;
				8'b1110000: c <= 9'b10110101;
				8'b1101001: c <= 9'b101000011;
				8'b1110011: c <= 9'b110111010;
				8'b1001100: c <= 9'b100010110;
				8'b100001: c <= 9'b1101010;
				8'b1000110: c <= 9'b111100001;
				8'b1110010: c <= 9'b1011;
				8'b1010000: c <= 9'b111111111;
				8'b1111010: c <= 9'b10110010;
				8'b1010101: c <= 9'b10110111;
				8'b111011: c <= 9'b11011011;
				8'b1001101: c <= 9'b10101001;
				8'b111111: c <= 9'b11110;
				8'b1101110: c <= 9'b10110111;
				8'b1111011: c <= 9'b11100000;
				8'b1001011: c <= 9'b110101110;
				8'b1101111: c <= 9'b100100101;
				8'b1101000: c <= 9'b100110111;
				8'b101100: c <= 9'b111111000;
				8'b100100: c <= 9'b110001000;
				8'b1111000: c <= 9'b101000;
				8'b1000101: c <= 9'b101011011;
				8'b1011001: c <= 9'b111100001;
				8'b110100: c <= 9'b101000110;
				8'b1111001: c <= 9'b11011100;
				8'b1110001: c <= 9'b11101011;
				8'b1001111: c <= 9'b111111111;
				8'b1100101: c <= 9'b11010001;
				8'b1111110: c <= 9'b1110111;
				8'b1111100: c <= 9'b101011101;
				8'b1010110: c <= 9'b101100100;
				8'b110010: c <= 9'b101000100;
				8'b1101101: c <= 9'b111011110;
				8'b100011: c <= 9'b101011110;
				8'b1110101: c <= 9'b10111010;
				8'b1111101: c <= 9'b111000101;
				8'b101001: c <= 9'b100010010;
				8'b1010010: c <= 9'b101000100;
				8'b1011000: c <= 9'b101100000;
				8'b101110: c <= 9'b11100110;
				8'b1000001: c <= 9'b110101001;
				default: c <= 9'b0;
			endcase
			9'b11011010 : case(di)
				8'b1000011: c <= 9'b1101001;
				8'b101000: c <= 9'b111010000;
				8'b111010: c <= 9'b101000011;
				8'b110110: c <= 9'b11111101;
				8'b1100100: c <= 9'b100001;
				8'b1000000: c <= 9'b11100010;
				8'b1110110: c <= 9'b111111101;
				8'b100101: c <= 9'b1100111;
				8'b101111: c <= 9'b11110;
				8'b100110: c <= 9'b110100101;
				8'b1100011: c <= 9'b101011001;
				8'b1001000: c <= 9'b111000010;
				8'b111000: c <= 9'b10010011;
				8'b110001: c <= 9'b10111111;
				8'b1010111: c <= 9'b10100100;
				8'b1001110: c <= 9'b10101001;
				8'b1101010: c <= 9'b11011000;
				8'b1001001: c <= 9'b110011100;
				8'b1100000: c <= 9'b111110001;
				8'b110111: c <= 9'b100010111;
				8'b1011101: c <= 9'b10101111;
				8'b1011011: c <= 9'b10011010;
				8'b111001: c <= 9'b101101;
				8'b1001010: c <= 9'b111101101;
				8'b110011: c <= 9'b111100101;
				8'b1101100: c <= 9'b101101000;
				8'b1110111: c <= 9'b100010110;
				8'b101011: c <= 9'b101100010;
				8'b1101011: c <= 9'b111111001;
				8'b111100: c <= 9'b110010;
				8'b1000111: c <= 9'b101000011;
				8'b1011111: c <= 9'b10101110;
				8'b1110100: c <= 9'b111011111;
				8'b101101: c <= 9'b110001100;
				8'b1010011: c <= 9'b101001001;
				8'b1100001: c <= 9'b111000111;
				8'b110101: c <= 9'b111111110;
				8'b1000100: c <= 9'b111010111;
				8'b1010001: c <= 9'b100010010;
				8'b1010100: c <= 9'b101011;
				8'b1100110: c <= 9'b10010000;
				8'b101010: c <= 9'b111000010;
				8'b1011110: c <= 9'b11001010;
				8'b1100111: c <= 9'b100010000;
				8'b1011010: c <= 9'b1001111;
				8'b1000010: c <= 9'b1100;
				8'b111101: c <= 9'b100101011;
				8'b110000: c <= 9'b11100011;
				8'b111110: c <= 9'b11001111;
				8'b1100010: c <= 9'b101100101;
				8'b1110000: c <= 9'b110111;
				8'b1101001: c <= 9'b110111111;
				8'b1110011: c <= 9'b110010101;
				8'b1001100: c <= 9'b110000010;
				8'b100001: c <= 9'b110111010;
				8'b1000110: c <= 9'b111000110;
				8'b1110010: c <= 9'b1110100;
				8'b1010000: c <= 9'b10001100;
				8'b1111010: c <= 9'b110001100;
				8'b1010101: c <= 9'b1010001;
				8'b111011: c <= 9'b1111000;
				8'b1001101: c <= 9'b10101;
				8'b111111: c <= 9'b110101100;
				8'b1101110: c <= 9'b110011101;
				8'b1111011: c <= 9'b11100110;
				8'b1001011: c <= 9'b101011111;
				8'b1101111: c <= 9'b110011010;
				8'b1101000: c <= 9'b1101010;
				8'b101100: c <= 9'b1010000;
				8'b100100: c <= 9'b111110101;
				8'b1111000: c <= 9'b111101010;
				8'b1000101: c <= 9'b100110111;
				8'b1011001: c <= 9'b111111110;
				8'b110100: c <= 9'b111110110;
				8'b1111001: c <= 9'b111111101;
				8'b1110001: c <= 9'b1011100;
				8'b1001111: c <= 9'b110011111;
				8'b1100101: c <= 9'b11001111;
				8'b1111110: c <= 9'b111100011;
				8'b1111100: c <= 9'b10011010;
				8'b1010110: c <= 9'b111100010;
				8'b110010: c <= 9'b11111010;
				8'b1101101: c <= 9'b100000111;
				8'b100011: c <= 9'b1110010;
				8'b1110101: c <= 9'b110010001;
				8'b1111101: c <= 9'b101010011;
				8'b101001: c <= 9'b111101001;
				8'b1010010: c <= 9'b10100111;
				8'b1011000: c <= 9'b10111011;
				8'b101110: c <= 9'b1001111;
				8'b1000001: c <= 9'b1011100;
				default: c <= 9'b0;
			endcase
			9'b110010 : case(di)
				8'b1000011: c <= 9'b1111000;
				8'b101000: c <= 9'b11111010;
				8'b111010: c <= 9'b11100100;
				8'b110110: c <= 9'b11001111;
				8'b1100100: c <= 9'b11000110;
				8'b1000000: c <= 9'b100101110;
				8'b1110110: c <= 9'b11010000;
				8'b100101: c <= 9'b111001111;
				8'b101111: c <= 9'b10111011;
				8'b100110: c <= 9'b100011010;
				8'b1100011: c <= 9'b110010101;
				8'b1001000: c <= 9'b10011010;
				8'b111000: c <= 9'b101001010;
				8'b110001: c <= 9'b1110100;
				8'b1010111: c <= 9'b110010010;
				8'b1001110: c <= 9'b11110111;
				8'b1101010: c <= 9'b10100111;
				8'b1001001: c <= 9'b1001100;
				8'b1100000: c <= 9'b100111010;
				8'b110111: c <= 9'b100100111;
				8'b1011101: c <= 9'b110000011;
				8'b1011011: c <= 9'b10111100;
				8'b111001: c <= 9'b100001010;
				8'b1001010: c <= 9'b111000011;
				8'b110011: c <= 9'b11010010;
				8'b1101100: c <= 9'b10111011;
				8'b1110111: c <= 9'b111110011;
				8'b101011: c <= 9'b11011110;
				8'b1101011: c <= 9'b10111010;
				8'b111100: c <= 9'b10000111;
				8'b1000111: c <= 9'b1111101;
				8'b1011111: c <= 9'b110010;
				8'b1110100: c <= 9'b111001000;
				8'b101101: c <= 9'b110010001;
				8'b1010011: c <= 9'b100101100;
				8'b1100001: c <= 9'b10101101;
				8'b110101: c <= 9'b100000010;
				8'b1000100: c <= 9'b11000010;
				8'b1010001: c <= 9'b101000110;
				8'b1010100: c <= 9'b11101011;
				8'b1100110: c <= 9'b100111011;
				8'b101010: c <= 9'b10011111;
				8'b1011110: c <= 9'b110100110;
				8'b1100111: c <= 9'b100100001;
				8'b1011010: c <= 9'b10010001;
				8'b1000010: c <= 9'b11110001;
				8'b111101: c <= 9'b10000001;
				8'b110000: c <= 9'b110101110;
				8'b111110: c <= 9'b11100101;
				8'b1100010: c <= 9'b100100000;
				8'b1110000: c <= 9'b101100111;
				8'b1101001: c <= 9'b10010110;
				8'b1110011: c <= 9'b111111011;
				8'b1001100: c <= 9'b10010000;
				8'b100001: c <= 9'b1110011;
				8'b1000110: c <= 9'b111110000;
				8'b1110010: c <= 9'b100101110;
				8'b1010000: c <= 9'b101111010;
				8'b1111010: c <= 9'b101000011;
				8'b1010101: c <= 9'b1100010;
				8'b111011: c <= 9'b110010001;
				8'b1001101: c <= 9'b10110001;
				8'b111111: c <= 9'b10000;
				8'b1101110: c <= 9'b110011010;
				8'b1111011: c <= 9'b110001;
				8'b1001011: c <= 9'b101000111;
				8'b1101111: c <= 9'b1100001;
				8'b1101000: c <= 9'b110101;
				8'b101100: c <= 9'b110010110;
				8'b100100: c <= 9'b10001000;
				8'b1111000: c <= 9'b110010100;
				8'b1000101: c <= 9'b101111001;
				8'b1011001: c <= 9'b10101000;
				8'b110100: c <= 9'b101011000;
				8'b1111001: c <= 9'b101111010;
				8'b1110001: c <= 9'b101100011;
				8'b1001111: c <= 9'b111010001;
				8'b1100101: c <= 9'b1111001;
				8'b1111110: c <= 9'b111101111;
				8'b1111100: c <= 9'b110111010;
				8'b1010110: c <= 9'b1100110;
				8'b110010: c <= 9'b111100000;
				8'b1101101: c <= 9'b110001101;
				8'b100011: c <= 9'b100100001;
				8'b1110101: c <= 9'b1011100;
				8'b1111101: c <= 9'b11001;
				8'b101001: c <= 9'b110010010;
				8'b1010010: c <= 9'b101100100;
				8'b1011000: c <= 9'b11101100;
				8'b101110: c <= 9'b101011111;
				8'b1000001: c <= 9'b111100001;
				default: c <= 9'b0;
			endcase
			9'b10010111 : case(di)
				8'b1000011: c <= 9'b101011111;
				8'b101000: c <= 9'b1110101;
				8'b111010: c <= 9'b100001100;
				8'b110110: c <= 9'b1010011;
				8'b1100100: c <= 9'b101101100;
				8'b1000000: c <= 9'b100000001;
				8'b1110110: c <= 9'b1110011;
				8'b100101: c <= 9'b111011001;
				8'b101111: c <= 9'b100011101;
				8'b100110: c <= 9'b100110011;
				8'b1100011: c <= 9'b101111010;
				8'b1001000: c <= 9'b11010001;
				8'b111000: c <= 9'b110010001;
				8'b110001: c <= 9'b110111011;
				8'b1010111: c <= 9'b110111;
				8'b1001110: c <= 9'b10000110;
				8'b1101010: c <= 9'b1111100;
				8'b1001001: c <= 9'b101101011;
				8'b1100000: c <= 9'b100110110;
				8'b110111: c <= 9'b11111;
				8'b1011101: c <= 9'b10101010;
				8'b1011011: c <= 9'b11100110;
				8'b111001: c <= 9'b101;
				8'b1001010: c <= 9'b111101001;
				8'b110011: c <= 9'b101110110;
				8'b1101100: c <= 9'b1110;
				8'b1110111: c <= 9'b10000;
				8'b101011: c <= 9'b100111010;
				8'b1101011: c <= 9'b10100000;
				8'b111100: c <= 9'b101;
				8'b1000111: c <= 9'b100101;
				8'b1011111: c <= 9'b110100011;
				8'b1110100: c <= 9'b111100101;
				8'b101101: c <= 9'b11111101;
				8'b1010011: c <= 9'b100100000;
				8'b1100001: c <= 9'b111001100;
				8'b110101: c <= 9'b110011100;
				8'b1000100: c <= 9'b101110010;
				8'b1010001: c <= 9'b111101100;
				8'b1010100: c <= 9'b101010001;
				8'b1100110: c <= 9'b11010010;
				8'b101010: c <= 9'b100101011;
				8'b1011110: c <= 9'b111100101;
				8'b1100111: c <= 9'b101110010;
				8'b1011010: c <= 9'b100100111;
				8'b1000010: c <= 9'b10010001;
				8'b111101: c <= 9'b110000001;
				8'b110000: c <= 9'b1101100;
				8'b111110: c <= 9'b101001100;
				8'b1100010: c <= 9'b10011000;
				8'b1110000: c <= 9'b100101100;
				8'b1101001: c <= 9'b100010100;
				8'b1110011: c <= 9'b110001000;
				8'b1001100: c <= 9'b10100;
				8'b100001: c <= 9'b11010;
				8'b1000110: c <= 9'b110111011;
				8'b1110010: c <= 9'b10010000;
				8'b1010000: c <= 9'b100111101;
				8'b1111010: c <= 9'b1001011;
				8'b1010101: c <= 9'b100010000;
				8'b111011: c <= 9'b101011001;
				8'b1001101: c <= 9'b111111001;
				8'b111111: c <= 9'b110100001;
				8'b1101110: c <= 9'b11111100;
				8'b1111011: c <= 9'b100100;
				8'b1001011: c <= 9'b101100110;
				8'b1101111: c <= 9'b11111000;
				8'b1101000: c <= 9'b111010001;
				8'b101100: c <= 9'b101000;
				8'b100100: c <= 9'b1010111;
				8'b1111000: c <= 9'b101010101;
				8'b1000101: c <= 9'b100101000;
				8'b1011001: c <= 9'b110110101;
				8'b110100: c <= 9'b111000110;
				8'b1111001: c <= 9'b110010;
				8'b1110001: c <= 9'b101001001;
				8'b1001111: c <= 9'b10000001;
				8'b1100101: c <= 9'b110011001;
				8'b1111110: c <= 9'b101001011;
				8'b1111100: c <= 9'b110010101;
				8'b1010110: c <= 9'b11010001;
				8'b110010: c <= 9'b100110101;
				8'b1101101: c <= 9'b111101010;
				8'b100011: c <= 9'b100110;
				8'b1110101: c <= 9'b1000;
				8'b1111101: c <= 9'b100101;
				8'b101001: c <= 9'b101001001;
				8'b1010010: c <= 9'b1101100;
				8'b1011000: c <= 9'b11000;
				8'b101110: c <= 9'b1111001;
				8'b1000001: c <= 9'b1111110;
				default: c <= 9'b0;
			endcase
			9'b1011110 : case(di)
				8'b1000011: c <= 9'b100010111;
				8'b101000: c <= 9'b111110110;
				8'b111010: c <= 9'b110011100;
				8'b110110: c <= 9'b1100100;
				8'b1100100: c <= 9'b111011110;
				8'b1000000: c <= 9'b1101;
				8'b1110110: c <= 9'b1100010;
				8'b100101: c <= 9'b110101;
				8'b101111: c <= 9'b100101110;
				8'b100110: c <= 9'b100010010;
				8'b1100011: c <= 9'b1101100;
				8'b1001000: c <= 9'b100001001;
				8'b111000: c <= 9'b10010100;
				8'b110001: c <= 9'b11000001;
				8'b1010111: c <= 9'b110001100;
				8'b1001110: c <= 9'b101011;
				8'b1101010: c <= 9'b111101100;
				8'b1001001: c <= 9'b110001001;
				8'b1100000: c <= 9'b101111111;
				8'b110111: c <= 9'b1110100;
				8'b1011101: c <= 9'b100111010;
				8'b1011011: c <= 9'b1110010;
				8'b111001: c <= 9'b11001000;
				8'b1001010: c <= 9'b100000111;
				8'b110011: c <= 9'b101001111;
				8'b1101100: c <= 9'b1111011;
				8'b1110111: c <= 9'b11001111;
				8'b101011: c <= 9'b111110000;
				8'b1101011: c <= 9'b100011011;
				8'b111100: c <= 9'b11001010;
				8'b1000111: c <= 9'b1001000;
				8'b1011111: c <= 9'b1001110;
				8'b1110100: c <= 9'b100110010;
				8'b101101: c <= 9'b111100000;
				8'b1010011: c <= 9'b11001000;
				8'b1100001: c <= 9'b11111100;
				8'b110101: c <= 9'b10000010;
				8'b1000100: c <= 9'b100001;
				8'b1010001: c <= 9'b10111;
				8'b1010100: c <= 9'b111111;
				8'b1100110: c <= 9'b101;
				8'b101010: c <= 9'b110100001;
				8'b1011110: c <= 9'b101110011;
				8'b1100111: c <= 9'b111110011;
				8'b1011010: c <= 9'b111000100;
				8'b1000010: c <= 9'b10101101;
				8'b111101: c <= 9'b101000010;
				8'b110000: c <= 9'b111010000;
				8'b111110: c <= 9'b11000111;
				8'b1100010: c <= 9'b1101111;
				8'b1110000: c <= 9'b100011011;
				8'b1101001: c <= 9'b11111000;
				8'b1110011: c <= 9'b11010001;
				8'b1001100: c <= 9'b11010010;
				8'b100001: c <= 9'b111010000;
				8'b1000110: c <= 9'b110000010;
				8'b1110010: c <= 9'b100001110;
				8'b1010000: c <= 9'b111011;
				8'b1111010: c <= 9'b100111001;
				8'b1010101: c <= 9'b10001001;
				8'b111011: c <= 9'b111000111;
				8'b1001101: c <= 9'b1111000;
				8'b111111: c <= 9'b10010111;
				8'b1101110: c <= 9'b101111010;
				8'b1111011: c <= 9'b110001101;
				8'b1001011: c <= 9'b11101000;
				8'b1101111: c <= 9'b11010010;
				8'b1101000: c <= 9'b111011011;
				8'b101100: c <= 9'b11101111;
				8'b100100: c <= 9'b1010010;
				8'b1111000: c <= 9'b110111011;
				8'b1000101: c <= 9'b110100001;
				8'b1011001: c <= 9'b110100001;
				8'b110100: c <= 9'b100010000;
				8'b1111001: c <= 9'b110101001;
				8'b1110001: c <= 9'b100011;
				8'b1001111: c <= 9'b1000;
				8'b1100101: c <= 9'b10010011;
				8'b1111110: c <= 9'b101011000;
				8'b1111100: c <= 9'b1100110;
				8'b1010110: c <= 9'b100010011;
				8'b110010: c <= 9'b101001000;
				8'b1101101: c <= 9'b11000000;
				8'b100011: c <= 9'b100101110;
				8'b1110101: c <= 9'b10101100;
				8'b1111101: c <= 9'b110011011;
				8'b101001: c <= 9'b11100011;
				8'b1010010: c <= 9'b111010000;
				8'b1011000: c <= 9'b11111;
				8'b101110: c <= 9'b110000110;
				8'b1000001: c <= 9'b100010001;
				default: c <= 9'b0;
			endcase
			9'b101010011 : case(di)
				8'b1000011: c <= 9'b10100000;
				8'b101000: c <= 9'b100000001;
				8'b111010: c <= 9'b10010011;
				8'b110110: c <= 9'b101001;
				8'b1100100: c <= 9'b100000011;
				8'b1000000: c <= 9'b11111011;
				8'b1110110: c <= 9'b11110010;
				8'b100101: c <= 9'b1111010;
				8'b101111: c <= 9'b10011100;
				8'b100110: c <= 9'b100101101;
				8'b1100011: c <= 9'b110001010;
				8'b1001000: c <= 9'b110111111;
				8'b111000: c <= 9'b111100011;
				8'b110001: c <= 9'b101110000;
				8'b1010111: c <= 9'b11100;
				8'b1001110: c <= 9'b101101110;
				8'b1101010: c <= 9'b11110111;
				8'b1001001: c <= 9'b101101011;
				8'b1100000: c <= 9'b1111101;
				8'b110111: c <= 9'b11100;
				8'b1011101: c <= 9'b111010010;
				8'b1011011: c <= 9'b100101;
				8'b111001: c <= 9'b101000111;
				8'b1001010: c <= 9'b11110011;
				8'b110011: c <= 9'b111000;
				8'b1101100: c <= 9'b110101111;
				8'b1110111: c <= 9'b111101110;
				8'b101011: c <= 9'b10100100;
				8'b1101011: c <= 9'b1100100;
				8'b111100: c <= 9'b111101110;
				8'b1000111: c <= 9'b1001101;
				8'b1011111: c <= 9'b11010;
				8'b1110100: c <= 9'b11101101;
				8'b101101: c <= 9'b101000100;
				8'b1010011: c <= 9'b111001011;
				8'b1100001: c <= 9'b100110100;
				8'b110101: c <= 9'b110000101;
				8'b1000100: c <= 9'b110100010;
				8'b1010001: c <= 9'b110100100;
				8'b1010100: c <= 9'b111100101;
				8'b1100110: c <= 9'b1111011;
				8'b101010: c <= 9'b11110;
				8'b1011110: c <= 9'b111001111;
				8'b1100111: c <= 9'b10111100;
				8'b1011010: c <= 9'b100110011;
				8'b1000010: c <= 9'b110011000;
				8'b111101: c <= 9'b100111111;
				8'b110000: c <= 9'b110100011;
				8'b111110: c <= 9'b101010111;
				8'b1100010: c <= 9'b111101110;
				8'b1110000: c <= 9'b11010101;
				8'b1101001: c <= 9'b101011011;
				8'b1110011: c <= 9'b1110101;
				8'b1001100: c <= 9'b101011101;
				8'b100001: c <= 9'b101001010;
				8'b1000110: c <= 9'b100011100;
				8'b1110010: c <= 9'b110011001;
				8'b1010000: c <= 9'b110010110;
				8'b1111010: c <= 9'b100001001;
				8'b1010101: c <= 9'b1010001;
				8'b111011: c <= 9'b111111000;
				8'b1001101: c <= 9'b101100010;
				8'b111111: c <= 9'b10011010;
				8'b1101110: c <= 9'b1101;
				8'b1111011: c <= 9'b111101;
				8'b1001011: c <= 9'b110111111;
				8'b1101111: c <= 9'b10100000;
				8'b1101000: c <= 9'b1100110;
				8'b101100: c <= 9'b11000;
				8'b100100: c <= 9'b11001010;
				8'b1111000: c <= 9'b110010101;
				8'b1000101: c <= 9'b11100010;
				8'b1011001: c <= 9'b10100110;
				8'b110100: c <= 9'b10101001;
				8'b1111001: c <= 9'b11110011;
				8'b1110001: c <= 9'b1111001;
				8'b1001111: c <= 9'b101001110;
				8'b1100101: c <= 9'b10110100;
				8'b1111110: c <= 9'b110111010;
				8'b1111100: c <= 9'b111101;
				8'b1010110: c <= 9'b101100;
				8'b110010: c <= 9'b100110011;
				8'b1101101: c <= 9'b110110010;
				8'b100011: c <= 9'b1000000;
				8'b1110101: c <= 9'b1111100;
				8'b1111101: c <= 9'b11000;
				8'b101001: c <= 9'b10111100;
				8'b1010010: c <= 9'b110010010;
				8'b1011000: c <= 9'b100101100;
				8'b101110: c <= 9'b110;
				8'b1000001: c <= 9'b10111010;
				default: c <= 9'b0;
			endcase
			9'b101101100 : case(di)
				8'b1000011: c <= 9'b100101011;
				8'b101000: c <= 9'b100110010;
				8'b111010: c <= 9'b10000000;
				8'b110110: c <= 9'b101011010;
				8'b1100100: c <= 9'b1100001;
				8'b1000000: c <= 9'b101111110;
				8'b1110110: c <= 9'b11110100;
				8'b100101: c <= 9'b10101;
				8'b101111: c <= 9'b10101001;
				8'b100110: c <= 9'b1100011;
				8'b1100011: c <= 9'b100011111;
				8'b1001000: c <= 9'b101111000;
				8'b111000: c <= 9'b100100010;
				8'b110001: c <= 9'b10101111;
				8'b1010111: c <= 9'b100101111;
				8'b1001110: c <= 9'b100111000;
				8'b1101010: c <= 9'b101011;
				8'b1001001: c <= 9'b1111111;
				8'b1100000: c <= 9'b101111000;
				8'b110111: c <= 9'b111101111;
				8'b1011101: c <= 9'b1100000;
				8'b1011011: c <= 9'b1;
				8'b111001: c <= 9'b101111010;
				8'b1001010: c <= 9'b100100;
				8'b110011: c <= 9'b11011000;
				8'b1101100: c <= 9'b11000001;
				8'b1110111: c <= 9'b101110110;
				8'b101011: c <= 9'b101101100;
				8'b1101011: c <= 9'b111010110;
				8'b111100: c <= 9'b111001111;
				8'b1000111: c <= 9'b101011000;
				8'b1011111: c <= 9'b10010011;
				8'b1110100: c <= 9'b100000010;
				8'b101101: c <= 9'b110001100;
				8'b1010011: c <= 9'b10011111;
				8'b1100001: c <= 9'b11011101;
				8'b110101: c <= 9'b11;
				8'b1000100: c <= 9'b100100001;
				8'b1010001: c <= 9'b11001011;
				8'b1010100: c <= 9'b11001010;
				8'b1100110: c <= 9'b10001100;
				8'b101010: c <= 9'b10001010;
				8'b1011110: c <= 9'b1011110;
				8'b1100111: c <= 9'b110011010;
				8'b1011010: c <= 9'b11100101;
				8'b1000010: c <= 9'b10111001;
				8'b111101: c <= 9'b110100001;
				8'b110000: c <= 9'b101101001;
				8'b111110: c <= 9'b10110111;
				8'b1100010: c <= 9'b111010100;
				8'b1110000: c <= 9'b101110111;
				8'b1101001: c <= 9'b110100100;
				8'b1110011: c <= 9'b11010010;
				8'b1001100: c <= 9'b100010110;
				8'b100001: c <= 9'b10001110;
				8'b1000110: c <= 9'b110011001;
				8'b1110010: c <= 9'b110011;
				8'b1010000: c <= 9'b10111100;
				8'b1111010: c <= 9'b10001010;
				8'b1010101: c <= 9'b111101111;
				8'b111011: c <= 9'b10111;
				8'b1001101: c <= 9'b111111111;
				8'b111111: c <= 9'b1110101;
				8'b1101110: c <= 9'b111100001;
				8'b1111011: c <= 9'b101011101;
				8'b1001011: c <= 9'b11001111;
				8'b1101111: c <= 9'b111111;
				8'b1101000: c <= 9'b110001100;
				8'b101100: c <= 9'b1100110;
				8'b100100: c <= 9'b100011100;
				8'b1111000: c <= 9'b100011010;
				8'b1000101: c <= 9'b10000011;
				8'b1011001: c <= 9'b111001100;
				8'b110100: c <= 9'b1110010;
				8'b1111001: c <= 9'b101001111;
				8'b1110001: c <= 9'b111101101;
				8'b1001111: c <= 9'b11111011;
				8'b1100101: c <= 9'b11001111;
				8'b1111110: c <= 9'b10010101;
				8'b1111100: c <= 9'b110110101;
				8'b1010110: c <= 9'b101011101;
				8'b110010: c <= 9'b1110111;
				8'b1101101: c <= 9'b110101010;
				8'b100011: c <= 9'b11111;
				8'b1110101: c <= 9'b111;
				8'b1111101: c <= 9'b101110111;
				8'b101001: c <= 9'b110100000;
				8'b1010010: c <= 9'b110010001;
				8'b1011000: c <= 9'b110;
				8'b101110: c <= 9'b111000100;
				8'b1000001: c <= 9'b10000111;
				default: c <= 9'b0;
			endcase
			9'b101101110 : case(di)
				8'b1000011: c <= 9'b100101101;
				8'b101000: c <= 9'b11001011;
				8'b111010: c <= 9'b100001011;
				8'b110110: c <= 9'b10110011;
				8'b1100100: c <= 9'b101010110;
				8'b1000000: c <= 9'b10011000;
				8'b1110110: c <= 9'b101101101;
				8'b100101: c <= 9'b100101100;
				8'b101111: c <= 9'b101;
				8'b100110: c <= 9'b1000100;
				8'b1100011: c <= 9'b111001010;
				8'b1001000: c <= 9'b100100010;
				8'b111000: c <= 9'b110101100;
				8'b110001: c <= 9'b11110000;
				8'b1010111: c <= 9'b110001;
				8'b1001110: c <= 9'b110110011;
				8'b1101010: c <= 9'b11010100;
				8'b1001001: c <= 9'b1111100;
				8'b1100000: c <= 9'b110000110;
				8'b110111: c <= 9'b100000100;
				8'b1011101: c <= 9'b111011011;
				8'b1011011: c <= 9'b100111110;
				8'b111001: c <= 9'b100010010;
				8'b1001010: c <= 9'b1001101;
				8'b110011: c <= 9'b111000101;
				8'b1101100: c <= 9'b10110010;
				8'b1110111: c <= 9'b1010010;
				8'b101011: c <= 9'b101011111;
				8'b1101011: c <= 9'b11111110;
				8'b111100: c <= 9'b11001101;
				8'b1000111: c <= 9'b110111011;
				8'b1011111: c <= 9'b1100110;
				8'b1110100: c <= 9'b101101010;
				8'b101101: c <= 9'b10001000;
				8'b1010011: c <= 9'b110010101;
				8'b1100001: c <= 9'b10000;
				8'b110101: c <= 9'b1101000;
				8'b1000100: c <= 9'b110001010;
				8'b1010001: c <= 9'b1110;
				8'b1010100: c <= 9'b101101100;
				8'b1100110: c <= 9'b110111001;
				8'b101010: c <= 9'b111000011;
				8'b1011110: c <= 9'b110000010;
				8'b1100111: c <= 9'b11111101;
				8'b1011010: c <= 9'b101110010;
				8'b1000010: c <= 9'b1010110;
				8'b111101: c <= 9'b10000000;
				8'b110000: c <= 9'b1011011;
				8'b111110: c <= 9'b10111001;
				8'b1100010: c <= 9'b100100111;
				8'b1110000: c <= 9'b10111101;
				8'b1101001: c <= 9'b1011110;
				8'b1110011: c <= 9'b1000;
				8'b1001100: c <= 9'b100;
				8'b100001: c <= 9'b100111111;
				8'b1000110: c <= 9'b1111100;
				8'b1110010: c <= 9'b101101;
				8'b1010000: c <= 9'b100111100;
				8'b1111010: c <= 9'b11101;
				8'b1010101: c <= 9'b1010001;
				8'b111011: c <= 9'b100110110;
				8'b1001101: c <= 9'b11100011;
				8'b111111: c <= 9'b100101001;
				8'b1101110: c <= 9'b110100110;
				8'b1111011: c <= 9'b111011;
				8'b1001011: c <= 9'b100100000;
				8'b1101111: c <= 9'b110110110;
				8'b1101000: c <= 9'b10011001;
				8'b101100: c <= 9'b100011101;
				8'b100100: c <= 9'b11111010;
				8'b1111000: c <= 9'b10001000;
				8'b1000101: c <= 9'b10000000;
				8'b1011001: c <= 9'b111011011;
				8'b110100: c <= 9'b110110011;
				8'b1111001: c <= 9'b100001100;
				8'b1110001: c <= 9'b110110;
				8'b1001111: c <= 9'b100101011;
				8'b1100101: c <= 9'b100111001;
				8'b1111110: c <= 9'b100110010;
				8'b1111100: c <= 9'b100100101;
				8'b1010110: c <= 9'b1101111;
				8'b110010: c <= 9'b10011001;
				8'b1101101: c <= 9'b11100;
				8'b100011: c <= 9'b100110111;
				8'b1110101: c <= 9'b111111;
				8'b1111101: c <= 9'b110001110;
				8'b101001: c <= 9'b110110;
				8'b1010010: c <= 9'b100011100;
				8'b1011000: c <= 9'b11110000;
				8'b101110: c <= 9'b10010111;
				8'b1000001: c <= 9'b110000101;
				default: c <= 9'b0;
			endcase
			9'b11001111 : case(di)
				8'b1000011: c <= 9'b10010100;
				8'b101000: c <= 9'b101001111;
				8'b111010: c <= 9'b101101110;
				8'b110110: c <= 9'b10100111;
				8'b1100100: c <= 9'b101000100;
				8'b1000000: c <= 9'b111001001;
				8'b1110110: c <= 9'b1011000;
				8'b100101: c <= 9'b110001110;
				8'b101111: c <= 9'b110011110;
				8'b100110: c <= 9'b111011110;
				8'b1100011: c <= 9'b100110100;
				8'b1001000: c <= 9'b11101011;
				8'b111000: c <= 9'b100010110;
				8'b110001: c <= 9'b110011111;
				8'b1010111: c <= 9'b101100001;
				8'b1001110: c <= 9'b111101;
				8'b1101010: c <= 9'b10111;
				8'b1001001: c <= 9'b101100010;
				8'b1100000: c <= 9'b11010001;
				8'b110111: c <= 9'b110111001;
				8'b1011101: c <= 9'b110010110;
				8'b1011011: c <= 9'b1100000;
				8'b111001: c <= 9'b1000101;
				8'b1001010: c <= 9'b1101100;
				8'b110011: c <= 9'b101101011;
				8'b1101100: c <= 9'b100011;
				8'b1110111: c <= 9'b1101;
				8'b101011: c <= 9'b101011101;
				8'b1101011: c <= 9'b101;
				8'b111100: c <= 9'b1100100;
				8'b1000111: c <= 9'b10010011;
				8'b1011111: c <= 9'b101010;
				8'b1110100: c <= 9'b110110111;
				8'b101101: c <= 9'b10000010;
				8'b1010011: c <= 9'b101100110;
				8'b1100001: c <= 9'b111010001;
				8'b110101: c <= 9'b101010100;
				8'b1000100: c <= 9'b111010010;
				8'b1010001: c <= 9'b110011000;
				8'b1010100: c <= 9'b1010111;
				8'b1100110: c <= 9'b111100000;
				8'b101010: c <= 9'b101001110;
				8'b1011110: c <= 9'b1100110;
				8'b1100111: c <= 9'b1100111;
				8'b1011010: c <= 9'b100101110;
				8'b1000010: c <= 9'b100001110;
				8'b111101: c <= 9'b10011101;
				8'b110000: c <= 9'b1000;
				8'b111110: c <= 9'b1010000;
				8'b1100010: c <= 9'b111100100;
				8'b1110000: c <= 9'b11;
				8'b1101001: c <= 9'b11011001;
				8'b1110011: c <= 9'b101110010;
				8'b1001100: c <= 9'b110101011;
				8'b100001: c <= 9'b110100111;
				8'b1000110: c <= 9'b100101100;
				8'b1110010: c <= 9'b1110111;
				8'b1010000: c <= 9'b1011;
				8'b1111010: c <= 9'b101001001;
				8'b1010101: c <= 9'b100111110;
				8'b111011: c <= 9'b101100100;
				8'b1001101: c <= 9'b101011110;
				8'b111111: c <= 9'b101111110;
				8'b1101110: c <= 9'b11001;
				8'b1111011: c <= 9'b11101011;
				8'b1001011: c <= 9'b101010010;
				8'b1101111: c <= 9'b11000;
				8'b1101000: c <= 9'b110101110;
				8'b101100: c <= 9'b10001001;
				8'b100100: c <= 9'b10001111;
				8'b1111000: c <= 9'b10101101;
				8'b1000101: c <= 9'b111100101;
				8'b1011001: c <= 9'b101011000;
				8'b110100: c <= 9'b100101110;
				8'b1111001: c <= 9'b110101101;
				8'b1110001: c <= 9'b1110011;
				8'b1001111: c <= 9'b11010100;
				8'b1100101: c <= 9'b100001010;
				8'b1111110: c <= 9'b101111110;
				8'b1111100: c <= 9'b11010001;
				8'b1010110: c <= 9'b100001010;
				8'b110010: c <= 9'b11000;
				8'b1101101: c <= 9'b1011110;
				8'b100011: c <= 9'b101100011;
				8'b1110101: c <= 9'b10001001;
				8'b1111101: c <= 9'b111100101;
				8'b101001: c <= 9'b101100110;
				8'b1010010: c <= 9'b100100010;
				8'b1011000: c <= 9'b111100010;
				8'b101110: c <= 9'b11000001;
				8'b1000001: c <= 9'b1010011;
				default: c <= 9'b0;
			endcase
			9'b101011101 : case(di)
				8'b1000011: c <= 9'b111010110;
				8'b101000: c <= 9'b1001101;
				8'b111010: c <= 9'b10111010;
				8'b110110: c <= 9'b111111001;
				8'b1100100: c <= 9'b100111001;
				8'b1000000: c <= 9'b11010000;
				8'b1110110: c <= 9'b100101011;
				8'b100101: c <= 9'b10100101;
				8'b101111: c <= 9'b1111100;
				8'b100110: c <= 9'b10010100;
				8'b1100011: c <= 9'b11110100;
				8'b1001000: c <= 9'b1101111;
				8'b111000: c <= 9'b100101100;
				8'b110001: c <= 9'b101100011;
				8'b1010111: c <= 9'b111000110;
				8'b1001110: c <= 9'b1111;
				8'b1101010: c <= 9'b11101101;
				8'b1001001: c <= 9'b1111000;
				8'b1100000: c <= 9'b111001111;
				8'b110111: c <= 9'b10001001;
				8'b1011101: c <= 9'b100001011;
				8'b1011011: c <= 9'b111000000;
				8'b111001: c <= 9'b10;
				8'b1001010: c <= 9'b11111001;
				8'b110011: c <= 9'b111110011;
				8'b1101100: c <= 9'b11100110;
				8'b1110111: c <= 9'b10110110;
				8'b101011: c <= 9'b101100101;
				8'b1101011: c <= 9'b10010110;
				8'b111100: c <= 9'b110000111;
				8'b1000111: c <= 9'b101001100;
				8'b1011111: c <= 9'b110010;
				8'b1110100: c <= 9'b101110000;
				8'b101101: c <= 9'b1111011;
				8'b1010011: c <= 9'b101101110;
				8'b1100001: c <= 9'b100001011;
				8'b110101: c <= 9'b10101;
				8'b1000100: c <= 9'b101011011;
				8'b1010001: c <= 9'b100110000;
				8'b1010100: c <= 9'b11100011;
				8'b1100110: c <= 9'b111110000;
				8'b101010: c <= 9'b111000100;
				8'b1011110: c <= 9'b101110011;
				8'b1100111: c <= 9'b101010101;
				8'b1011010: c <= 9'b11001;
				8'b1000010: c <= 9'b101110010;
				8'b111101: c <= 9'b110100100;
				8'b110000: c <= 9'b111101111;
				8'b111110: c <= 9'b111000010;
				8'b1100010: c <= 9'b111111111;
				8'b1110000: c <= 9'b1100100;
				8'b1101001: c <= 9'b1011011;
				8'b1110011: c <= 9'b1011111;
				8'b1001100: c <= 9'b10001011;
				8'b100001: c <= 9'b10111101;
				8'b1000110: c <= 9'b110110;
				8'b1110010: c <= 9'b1010001;
				8'b1010000: c <= 9'b111010010;
				8'b1111010: c <= 9'b10011;
				8'b1010101: c <= 9'b100000010;
				8'b111011: c <= 9'b11001010;
				8'b1001101: c <= 9'b111001011;
				8'b111111: c <= 9'b111110001;
				8'b1101110: c <= 9'b101011101;
				8'b1111011: c <= 9'b1100;
				8'b1001011: c <= 9'b11110110;
				8'b1101111: c <= 9'b110111100;
				8'b1101000: c <= 9'b110011100;
				8'b101100: c <= 9'b110101100;
				8'b100100: c <= 9'b11101001;
				8'b1111000: c <= 9'b100101011;
				8'b1000101: c <= 9'b100010110;
				8'b1011001: c <= 9'b100110100;
				8'b110100: c <= 9'b1001010;
				8'b1111001: c <= 9'b111000100;
				8'b1110001: c <= 9'b101101;
				8'b1001111: c <= 9'b110001110;
				8'b1100101: c <= 9'b111001001;
				8'b1111110: c <= 9'b100011001;
				8'b1111100: c <= 9'b110111111;
				8'b1010110: c <= 9'b100000001;
				8'b110010: c <= 9'b101010001;
				8'b1101101: c <= 9'b100100110;
				8'b100011: c <= 9'b111000010;
				8'b1110101: c <= 9'b1011011;
				8'b1111101: c <= 9'b11011000;
				8'b101001: c <= 9'b110001100;
				8'b1010010: c <= 9'b101001011;
				8'b1011000: c <= 9'b111111110;
				8'b101110: c <= 9'b11011010;
				8'b1000001: c <= 9'b110000000;
				default: c <= 9'b0;
			endcase
			9'b110111110 : case(di)
				8'b1000011: c <= 9'b110010010;
				8'b101000: c <= 9'b1111001;
				8'b111010: c <= 9'b100010101;
				8'b110110: c <= 9'b101110000;
				8'b1100100: c <= 9'b1101001;
				8'b1000000: c <= 9'b11111000;
				8'b1110110: c <= 9'b1011110;
				8'b100101: c <= 9'b11111010;
				8'b101111: c <= 9'b1011010;
				8'b100110: c <= 9'b10110101;
				8'b1100011: c <= 9'b110100100;
				8'b1001000: c <= 9'b10111001;
				8'b111000: c <= 9'b111001001;
				8'b110001: c <= 9'b10010000;
				8'b1010111: c <= 9'b10101101;
				8'b1001110: c <= 9'b110110000;
				8'b1101010: c <= 9'b10101100;
				8'b1001001: c <= 9'b100010100;
				8'b1100000: c <= 9'b10100100;
				8'b110111: c <= 9'b111000011;
				8'b1011101: c <= 9'b101001111;
				8'b1011011: c <= 9'b100110;
				8'b111001: c <= 9'b100111000;
				8'b1001010: c <= 9'b101101000;
				8'b110011: c <= 9'b1100001;
				8'b1101100: c <= 9'b1110010;
				8'b1110111: c <= 9'b100010;
				8'b101011: c <= 9'b100100001;
				8'b1101011: c <= 9'b100101;
				8'b111100: c <= 9'b110110111;
				8'b1000111: c <= 9'b100111001;
				8'b1011111: c <= 9'b10001110;
				8'b1110100: c <= 9'b111111000;
				8'b101101: c <= 9'b11111110;
				8'b1010011: c <= 9'b100010010;
				8'b1100001: c <= 9'b111100100;
				8'b110101: c <= 9'b10111000;
				8'b1000100: c <= 9'b10110001;
				8'b1010001: c <= 9'b100000111;
				8'b1010100: c <= 9'b11110010;
				8'b1100110: c <= 9'b111001110;
				8'b101010: c <= 9'b100;
				8'b1011110: c <= 9'b10101011;
				8'b1100111: c <= 9'b10111100;
				8'b1011010: c <= 9'b10101011;
				8'b1000010: c <= 9'b101001011;
				8'b111101: c <= 9'b100001001;
				8'b110000: c <= 9'b100111101;
				8'b111110: c <= 9'b1010000;
				8'b1100010: c <= 9'b111110000;
				8'b1110000: c <= 9'b101010001;
				8'b1101001: c <= 9'b101100111;
				8'b1110011: c <= 9'b11111110;
				8'b1001100: c <= 9'b101011001;
				8'b100001: c <= 9'b10000111;
				8'b1000110: c <= 9'b1010101;
				8'b1110010: c <= 9'b11011001;
				8'b1010000: c <= 9'b100011100;
				8'b1111010: c <= 9'b101001110;
				8'b1010101: c <= 9'b110101001;
				8'b111011: c <= 9'b101011111;
				8'b1001101: c <= 9'b11011001;
				8'b111111: c <= 9'b11010101;
				8'b1101110: c <= 9'b100110110;
				8'b1111011: c <= 9'b1110;
				8'b1001011: c <= 9'b1010011;
				8'b1101111: c <= 9'b10100100;
				8'b1101000: c <= 9'b10101;
				8'b101100: c <= 9'b111011011;
				8'b100100: c <= 9'b111000010;
				8'b1111000: c <= 9'b110001010;
				8'b1000101: c <= 9'b101000110;
				8'b1011001: c <= 9'b101010010;
				8'b110100: c <= 9'b110100101;
				8'b1111001: c <= 9'b101101001;
				8'b1110001: c <= 9'b1011111;
				8'b1001111: c <= 9'b100000110;
				8'b1100101: c <= 9'b1101110;
				8'b1111110: c <= 9'b1000;
				8'b1111100: c <= 9'b101001000;
				8'b1010110: c <= 9'b111111;
				8'b110010: c <= 9'b1111011;
				8'b1101101: c <= 9'b10111001;
				8'b100011: c <= 9'b1001;
				8'b1110101: c <= 9'b101110101;
				8'b1111101: c <= 9'b110111111;
				8'b101001: c <= 9'b1001001;
				8'b1010010: c <= 9'b10001111;
				8'b1011000: c <= 9'b1001001;
				8'b101110: c <= 9'b111111101;
				8'b1000001: c <= 9'b1000001;
				default: c <= 9'b0;
			endcase
			9'b101001000 : case(di)
				8'b1000011: c <= 9'b1110111;
				8'b101000: c <= 9'b10010101;
				8'b111010: c <= 9'b100110110;
				8'b110110: c <= 9'b111101100;
				8'b1100100: c <= 9'b101011;
				8'b1000000: c <= 9'b110011110;
				8'b1110110: c <= 9'b10111110;
				8'b100101: c <= 9'b111100000;
				8'b101111: c <= 9'b10110;
				8'b100110: c <= 9'b111100010;
				8'b1100011: c <= 9'b11110000;
				8'b1001000: c <= 9'b100101110;
				8'b111000: c <= 9'b1100001;
				8'b110001: c <= 9'b1110000;
				8'b1010111: c <= 9'b1001110;
				8'b1001110: c <= 9'b1000011;
				8'b1101010: c <= 9'b110111111;
				8'b1001001: c <= 9'b10001101;
				8'b1100000: c <= 9'b111010100;
				8'b110111: c <= 9'b110010010;
				8'b1011101: c <= 9'b110011101;
				8'b1011011: c <= 9'b1001000;
				8'b111001: c <= 9'b11100011;
				8'b1001010: c <= 9'b11010101;
				8'b110011: c <= 9'b11100010;
				8'b1101100: c <= 9'b101110101;
				8'b1110111: c <= 9'b11111100;
				8'b101011: c <= 9'b1101110;
				8'b1101011: c <= 9'b101100110;
				8'b111100: c <= 9'b110010101;
				8'b1000111: c <= 9'b10011;
				8'b1011111: c <= 9'b111011010;
				8'b1110100: c <= 9'b110010100;
				8'b101101: c <= 9'b101110101;
				8'b1010011: c <= 9'b100000111;
				8'b1100001: c <= 9'b110000010;
				8'b110101: c <= 9'b11100011;
				8'b1000100: c <= 9'b110001011;
				8'b1010001: c <= 9'b100111011;
				8'b1010100: c <= 9'b111100100;
				8'b1100110: c <= 9'b110111;
				8'b101010: c <= 9'b10010;
				8'b1011110: c <= 9'b10100100;
				8'b1100111: c <= 9'b1101010;
				8'b1011010: c <= 9'b101000010;
				8'b1000010: c <= 9'b10101000;
				8'b111101: c <= 9'b101110000;
				8'b110000: c <= 9'b1110111;
				8'b111110: c <= 9'b101011;
				8'b1100010: c <= 9'b100000000;
				8'b1110000: c <= 9'b10011000;
				8'b1101001: c <= 9'b101111110;
				8'b1110011: c <= 9'b10001011;
				8'b1001100: c <= 9'b110100011;
				8'b100001: c <= 9'b110001111;
				8'b1000110: c <= 9'b110010011;
				8'b1110010: c <= 9'b111010111;
				8'b1010000: c <= 9'b11011000;
				8'b1111010: c <= 9'b10000001;
				8'b1010101: c <= 9'b101011001;
				8'b111011: c <= 9'b10011;
				8'b1001101: c <= 9'b100010001;
				8'b111111: c <= 9'b11011110;
				8'b1101110: c <= 9'b11011110;
				8'b1111011: c <= 9'b101001;
				8'b1001011: c <= 9'b110110101;
				8'b1101111: c <= 9'b11111000;
				8'b1101000: c <= 9'b101111110;
				8'b101100: c <= 9'b1011010;
				8'b100100: c <= 9'b111001011;
				8'b1111000: c <= 9'b10111;
				8'b1000101: c <= 9'b111001011;
				8'b1011001: c <= 9'b10111100;
				8'b110100: c <= 9'b110001110;
				8'b1111001: c <= 9'b110101101;
				8'b1110001: c <= 9'b10010001;
				8'b1001111: c <= 9'b1011100;
				8'b1100101: c <= 9'b11001110;
				8'b1111110: c <= 9'b101110101;
				8'b1111100: c <= 9'b11000111;
				8'b1010110: c <= 9'b10100;
				8'b110010: c <= 9'b10101110;
				8'b1101101: c <= 9'b1011000;
				8'b100011: c <= 9'b110011000;
				8'b1110101: c <= 9'b11011010;
				8'b1111101: c <= 9'b100001011;
				8'b101001: c <= 9'b11101000;
				8'b1010010: c <= 9'b110010110;
				8'b1011000: c <= 9'b110001100;
				8'b101110: c <= 9'b11011;
				8'b1000001: c <= 9'b11001100;
				default: c <= 9'b0;
			endcase
			9'b100010111 : case(di)
				8'b1000011: c <= 9'b11001100;
				8'b101000: c <= 9'b1111011;
				8'b111010: c <= 9'b111000100;
				8'b110110: c <= 9'b1101100;
				8'b1100100: c <= 9'b100001100;
				8'b1000000: c <= 9'b11100;
				8'b1110110: c <= 9'b1000011;
				8'b100101: c <= 9'b10101110;
				8'b101111: c <= 9'b1110001;
				8'b100110: c <= 9'b100111010;
				8'b1100011: c <= 9'b11111011;
				8'b1001000: c <= 9'b110010111;
				8'b111000: c <= 9'b110101010;
				8'b110001: c <= 9'b111010110;
				8'b1010111: c <= 9'b101010110;
				8'b1001110: c <= 9'b10001010;
				8'b1101010: c <= 9'b111101;
				8'b1001001: c <= 9'b10011100;
				8'b1100000: c <= 9'b111101;
				8'b110111: c <= 9'b101010001;
				8'b1011101: c <= 9'b110110100;
				8'b1011011: c <= 9'b111001000;
				8'b111001: c <= 9'b101010001;
				8'b1001010: c <= 9'b10010111;
				8'b110011: c <= 9'b111000110;
				8'b1101100: c <= 9'b1100111;
				8'b1110111: c <= 9'b101100000;
				8'b101011: c <= 9'b1100110;
				8'b1101011: c <= 9'b110111;
				8'b111100: c <= 9'b111101;
				8'b1000111: c <= 9'b1010010;
				8'b1011111: c <= 9'b1000010;
				8'b1110100: c <= 9'b111010100;
				8'b101101: c <= 9'b111001;
				8'b1010011: c <= 9'b111110000;
				8'b1100001: c <= 9'b10111110;
				8'b110101: c <= 9'b1001001;
				8'b1000100: c <= 9'b111101110;
				8'b1010001: c <= 9'b110100;
				8'b1010100: c <= 9'b111000000;
				8'b1100110: c <= 9'b110011100;
				8'b101010: c <= 9'b111010110;
				8'b1011110: c <= 9'b10110001;
				8'b1100111: c <= 9'b100000101;
				8'b1011010: c <= 9'b110111100;
				8'b1000010: c <= 9'b111010001;
				8'b111101: c <= 9'b110001000;
				8'b110000: c <= 9'b110011111;
				8'b111110: c <= 9'b10100101;
				8'b1100010: c <= 9'b111101110;
				8'b1110000: c <= 9'b100010000;
				8'b1101001: c <= 9'b111111111;
				8'b1110011: c <= 9'b1101001;
				8'b1001100: c <= 9'b11011000;
				8'b100001: c <= 9'b111111101;
				8'b1000110: c <= 9'b10110;
				8'b1110010: c <= 9'b111100011;
				8'b1010000: c <= 9'b101001;
				8'b1111010: c <= 9'b110110010;
				8'b1010101: c <= 9'b1000100;
				8'b111011: c <= 9'b111001010;
				8'b1001101: c <= 9'b10010000;
				8'b111111: c <= 9'b10001100;
				8'b1101110: c <= 9'b11011011;
				8'b1111011: c <= 9'b10000010;
				8'b1001011: c <= 9'b1011110;
				8'b1101111: c <= 9'b10101010;
				8'b1101000: c <= 9'b110010100;
				8'b101100: c <= 9'b100000011;
				8'b100100: c <= 9'b101101001;
				8'b1111000: c <= 9'b111110001;
				8'b1000101: c <= 9'b110101010;
				8'b1011001: c <= 9'b1110001;
				8'b110100: c <= 9'b111111;
				8'b1111001: c <= 9'b10001101;
				8'b1110001: c <= 9'b110111000;
				8'b1001111: c <= 9'b100011000;
				8'b1100101: c <= 9'b100111111;
				8'b1111110: c <= 9'b100111010;
				8'b1111100: c <= 9'b110100;
				8'b1010110: c <= 9'b110100110;
				8'b110010: c <= 9'b11100111;
				8'b1101101: c <= 9'b110101011;
				8'b100011: c <= 9'b101000101;
				8'b1110101: c <= 9'b110100;
				8'b1111101: c <= 9'b10011001;
				8'b101001: c <= 9'b10100111;
				8'b1010010: c <= 9'b101111110;
				8'b1011000: c <= 9'b100110000;
				8'b101110: c <= 9'b101110011;
				8'b1000001: c <= 9'b110100100;
				default: c <= 9'b0;
			endcase
			9'b101111110 : case(di)
				8'b1000011: c <= 9'b110110011;
				8'b101000: c <= 9'b1100101;
				8'b111010: c <= 9'b100000111;
				8'b110110: c <= 9'b10000000;
				8'b1100100: c <= 9'b10110100;
				8'b1000000: c <= 9'b11110110;
				8'b1110110: c <= 9'b110011;
				8'b100101: c <= 9'b101010010;
				8'b101111: c <= 9'b101100101;
				8'b100110: c <= 9'b110010111;
				8'b1100011: c <= 9'b101;
				8'b1001000: c <= 9'b110001111;
				8'b111000: c <= 9'b1101000;
				8'b110001: c <= 9'b11100111;
				8'b1010111: c <= 9'b101101000;
				8'b1001110: c <= 9'b111111101;
				8'b1101010: c <= 9'b10100111;
				8'b1001001: c <= 9'b100100010;
				8'b1100000: c <= 9'b110100111;
				8'b110111: c <= 9'b10010011;
				8'b1011101: c <= 9'b110110110;
				8'b1011011: c <= 9'b1010001;
				8'b111001: c <= 9'b100000001;
				8'b1001010: c <= 9'b11000100;
				8'b110011: c <= 9'b100110110;
				8'b1101100: c <= 9'b100110111;
				8'b1110111: c <= 9'b111000000;
				8'b101011: c <= 9'b100100;
				8'b1101011: c <= 9'b100000101;
				8'b111100: c <= 9'b1010001;
				8'b1000111: c <= 9'b100000011;
				8'b1011111: c <= 9'b110101010;
				8'b1110100: c <= 9'b10111110;
				8'b101101: c <= 9'b11010111;
				8'b1010011: c <= 9'b111000110;
				8'b1100001: c <= 9'b110000101;
				8'b110101: c <= 9'b111011011;
				8'b1000100: c <= 9'b101001111;
				8'b1010001: c <= 9'b11111011;
				8'b1010100: c <= 9'b110101110;
				8'b1100110: c <= 9'b110001;
				8'b101010: c <= 9'b11111011;
				8'b1011110: c <= 9'b11010101;
				8'b1100111: c <= 9'b11111001;
				8'b1011010: c <= 9'b101011000;
				8'b1000010: c <= 9'b111011100;
				8'b111101: c <= 9'b1010001;
				8'b110000: c <= 9'b110011100;
				8'b111110: c <= 9'b10000001;
				8'b1100010: c <= 9'b101000110;
				8'b1110000: c <= 9'b100101011;
				8'b1101001: c <= 9'b111010;
				8'b1110011: c <= 9'b101000101;
				8'b1001100: c <= 9'b11100010;
				8'b100001: c <= 9'b110100111;
				8'b1000110: c <= 9'b1111110;
				8'b1110010: c <= 9'b1101;
				8'b1010000: c <= 9'b101100101;
				8'b1111010: c <= 9'b11011;
				8'b1010101: c <= 9'b100110000;
				8'b111011: c <= 9'b110000001;
				8'b1001101: c <= 9'b1100111;
				8'b111111: c <= 9'b110100;
				8'b1101110: c <= 9'b10111;
				8'b1111011: c <= 9'b100100001;
				8'b1001011: c <= 9'b110011000;
				8'b1101111: c <= 9'b11110111;
				8'b1101000: c <= 9'b110001110;
				8'b101100: c <= 9'b111110000;
				8'b100100: c <= 9'b111100001;
				8'b1111000: c <= 9'b1101001;
				8'b1000101: c <= 9'b101101;
				8'b1011001: c <= 9'b111011111;
				8'b110100: c <= 9'b111001000;
				8'b1111001: c <= 9'b11011001;
				8'b1110001: c <= 9'b110101010;
				8'b1001111: c <= 9'b10011111;
				8'b1100101: c <= 9'b110001111;
				8'b1111110: c <= 9'b1110100;
				8'b1111100: c <= 9'b11010011;
				8'b1010110: c <= 9'b11100111;
				8'b110010: c <= 9'b100111111;
				8'b1101101: c <= 9'b101101100;
				8'b100011: c <= 9'b111001010;
				8'b1110101: c <= 9'b1000010;
				8'b1111101: c <= 9'b110000000;
				8'b101001: c <= 9'b101101001;
				8'b1010010: c <= 9'b110010001;
				8'b1011000: c <= 9'b111000011;
				8'b101110: c <= 9'b101000110;
				8'b1000001: c <= 9'b110001100;
				default: c <= 9'b0;
			endcase
			9'b11000111 : case(di)
				8'b1000011: c <= 9'b101001000;
				8'b101000: c <= 9'b100000101;
				8'b111010: c <= 9'b100011101;
				8'b110110: c <= 9'b111001001;
				8'b1100100: c <= 9'b110001;
				8'b1000000: c <= 9'b1111010;
				8'b1110110: c <= 9'b11010111;
				8'b100101: c <= 9'b101111001;
				8'b101111: c <= 9'b111000101;
				8'b100110: c <= 9'b11101111;
				8'b1100011: c <= 9'b110000010;
				8'b1001000: c <= 9'b1101110;
				8'b111000: c <= 9'b100011;
				8'b110001: c <= 9'b110110010;
				8'b1010111: c <= 9'b111010;
				8'b1001110: c <= 9'b110110111;
				8'b1101010: c <= 9'b11101100;
				8'b1001001: c <= 9'b101100010;
				8'b1100000: c <= 9'b11011011;
				8'b110111: c <= 9'b110011011;
				8'b1011101: c <= 9'b1110101;
				8'b1011011: c <= 9'b101111110;
				8'b111001: c <= 9'b10011010;
				8'b1001010: c <= 9'b1000011;
				8'b110011: c <= 9'b100000000;
				8'b1101100: c <= 9'b10111;
				8'b1110111: c <= 9'b10101101;
				8'b101011: c <= 9'b111110011;
				8'b1101011: c <= 9'b11000001;
				8'b111100: c <= 9'b100011111;
				8'b1000111: c <= 9'b10101110;
				8'b1011111: c <= 9'b111011001;
				8'b1110100: c <= 9'b1110011;
				8'b101101: c <= 9'b101000111;
				8'b1010011: c <= 9'b10101000;
				8'b1100001: c <= 9'b101101110;
				8'b110101: c <= 9'b110001;
				8'b1000100: c <= 9'b101011011;
				8'b1010001: c <= 9'b110010110;
				8'b1010100: c <= 9'b110100001;
				8'b1100110: c <= 9'b100100110;
				8'b101010: c <= 9'b1000001;
				8'b1011110: c <= 9'b110001011;
				8'b1100111: c <= 9'b11101000;
				8'b1011010: c <= 9'b111111101;
				8'b1000010: c <= 9'b111101001;
				8'b111101: c <= 9'b111100111;
				8'b110000: c <= 9'b11111100;
				8'b111110: c <= 9'b100000100;
				8'b1100010: c <= 9'b1111100;
				8'b1110000: c <= 9'b110011;
				8'b1101001: c <= 9'b1000010;
				8'b1110011: c <= 9'b11010100;
				8'b1001100: c <= 9'b11111010;
				8'b100001: c <= 9'b111100110;
				8'b1000110: c <= 9'b1111101;
				8'b1110010: c <= 9'b101000111;
				8'b1010000: c <= 9'b100110101;
				8'b1111010: c <= 9'b100111111;
				8'b1010101: c <= 9'b110111100;
				8'b111011: c <= 9'b101010111;
				8'b1001101: c <= 9'b1001100;
				8'b111111: c <= 9'b1001;
				8'b1101110: c <= 9'b10111110;
				8'b1111011: c <= 9'b100111110;
				8'b1001011: c <= 9'b111001101;
				8'b1101111: c <= 9'b1000100;
				8'b1101000: c <= 9'b111011100;
				8'b101100: c <= 9'b100001;
				8'b100100: c <= 9'b10101010;
				8'b1111000: c <= 9'b100010110;
				8'b1000101: c <= 9'b11001101;
				8'b1011001: c <= 9'b110001111;
				8'b110100: c <= 9'b1000000;
				8'b1111001: c <= 9'b100010100;
				8'b1110001: c <= 9'b101100110;
				8'b1001111: c <= 9'b11011000;
				8'b1100101: c <= 9'b10001010;
				8'b1111110: c <= 9'b100010110;
				8'b1111100: c <= 9'b10000101;
				8'b1010110: c <= 9'b111110000;
				8'b110010: c <= 9'b1110011;
				8'b1101101: c <= 9'b110111110;
				8'b100011: c <= 9'b1000000;
				8'b1110101: c <= 9'b110001000;
				8'b1111101: c <= 9'b110000111;
				8'b101001: c <= 9'b101100010;
				8'b1010010: c <= 9'b100101000;
				8'b1011000: c <= 9'b101000;
				8'b101110: c <= 9'b101001001;
				8'b1000001: c <= 9'b100100001;
				default: c <= 9'b0;
			endcase
			9'b10111000 : case(di)
				8'b1000011: c <= 9'b101110111;
				8'b101000: c <= 9'b1110100;
				8'b111010: c <= 9'b11010111;
				8'b110110: c <= 9'b110111110;
				8'b1100100: c <= 9'b100100000;
				8'b1000000: c <= 9'b11111000;
				8'b1110110: c <= 9'b111111000;
				8'b100101: c <= 9'b100011000;
				8'b101111: c <= 9'b111101010;
				8'b100110: c <= 9'b110100010;
				8'b1100011: c <= 9'b100100111;
				8'b1001000: c <= 9'b101001000;
				8'b111000: c <= 9'b110010111;
				8'b110001: c <= 9'b101011111;
				8'b1010111: c <= 9'b10001100;
				8'b1001110: c <= 9'b10110110;
				8'b1101010: c <= 9'b10100101;
				8'b1001001: c <= 9'b11110001;
				8'b1100000: c <= 9'b100001010;
				8'b110111: c <= 9'b100101100;
				8'b1011101: c <= 9'b11111001;
				8'b1011011: c <= 9'b111011111;
				8'b111001: c <= 9'b1011011;
				8'b1001010: c <= 9'b1;
				8'b110011: c <= 9'b1001000;
				8'b1101100: c <= 9'b101001100;
				8'b1110111: c <= 9'b10001110;
				8'b101011: c <= 9'b111100111;
				8'b1101011: c <= 9'b101001110;
				8'b111100: c <= 9'b110010010;
				8'b1000111: c <= 9'b10101110;
				8'b1011111: c <= 9'b111111011;
				8'b1110100: c <= 9'b101100011;
				8'b101101: c <= 9'b110010110;
				8'b1010011: c <= 9'b101101011;
				8'b1100001: c <= 9'b1010110;
				8'b110101: c <= 9'b101001;
				8'b1000100: c <= 9'b1111111;
				8'b1010001: c <= 9'b10000011;
				8'b1010100: c <= 9'b111110001;
				8'b1100110: c <= 9'b11100;
				8'b101010: c <= 9'b1000010;
				8'b1011110: c <= 9'b110000101;
				8'b1100111: c <= 9'b100110010;
				8'b1011010: c <= 9'b110010001;
				8'b1000010: c <= 9'b111000111;
				8'b111101: c <= 9'b1111011;
				8'b110000: c <= 9'b11001010;
				8'b111110: c <= 9'b101001011;
				8'b1100010: c <= 9'b1100110;
				8'b1110000: c <= 9'b101110000;
				8'b1101001: c <= 9'b1111100;
				8'b1110011: c <= 9'b10001001;
				8'b1001100: c <= 9'b10111001;
				8'b100001: c <= 9'b100111011;
				8'b1000110: c <= 9'b110100010;
				8'b1110010: c <= 9'b100001101;
				8'b1010000: c <= 9'b101001111;
				8'b1111010: c <= 9'b110100;
				8'b1010101: c <= 9'b110010110;
				8'b111011: c <= 9'b111110000;
				8'b1001101: c <= 9'b111100101;
				8'b111111: c <= 9'b110011000;
				8'b1101110: c <= 9'b1111011;
				8'b1111011: c <= 9'b100100011;
				8'b1001011: c <= 9'b111111010;
				8'b1101111: c <= 9'b101010101;
				8'b1101000: c <= 9'b111101001;
				8'b101100: c <= 9'b11000001;
				8'b100100: c <= 9'b11110011;
				8'b1111000: c <= 9'b10010;
				8'b1000101: c <= 9'b110011100;
				8'b1011001: c <= 9'b110110110;
				8'b110100: c <= 9'b110001110;
				8'b1111001: c <= 9'b10001011;
				8'b1110001: c <= 9'b110011110;
				8'b1001111: c <= 9'b111101100;
				8'b1100101: c <= 9'b111001000;
				8'b1111110: c <= 9'b111011001;
				8'b1111100: c <= 9'b1001111;
				8'b1010110: c <= 9'b111011011;
				8'b110010: c <= 9'b101100001;
				8'b1101101: c <= 9'b100011101;
				8'b100011: c <= 9'b101110001;
				8'b1110101: c <= 9'b100011101;
				8'b1111101: c <= 9'b100100;
				8'b101001: c <= 9'b11000011;
				8'b1010010: c <= 9'b110101110;
				8'b1011000: c <= 9'b111011;
				8'b101110: c <= 9'b101111000;
				8'b1000001: c <= 9'b110111001;
				default: c <= 9'b0;
			endcase
			9'b110101110 : case(di)
				8'b1000011: c <= 9'b11100101;
				8'b101000: c <= 9'b101101110;
				8'b111010: c <= 9'b110011110;
				8'b110110: c <= 9'b111010110;
				8'b1100100: c <= 9'b100100110;
				8'b1000000: c <= 9'b11100011;
				8'b1110110: c <= 9'b110011000;
				8'b100101: c <= 9'b10000001;
				8'b101111: c <= 9'b111101111;
				8'b100110: c <= 9'b111000011;
				8'b1100011: c <= 9'b1011011;
				8'b1001000: c <= 9'b110011111;
				8'b111000: c <= 9'b111010110;
				8'b110001: c <= 9'b101100;
				8'b1010111: c <= 9'b101001011;
				8'b1001110: c <= 9'b10110101;
				8'b1101010: c <= 9'b1001111;
				8'b1001001: c <= 9'b111110101;
				8'b1100000: c <= 9'b1111000;
				8'b110111: c <= 9'b111111101;
				8'b1011101: c <= 9'b100001100;
				8'b1011011: c <= 9'b1000;
				8'b111001: c <= 9'b100011000;
				8'b1001010: c <= 9'b101100000;
				8'b110011: c <= 9'b111100011;
				8'b1101100: c <= 9'b110100001;
				8'b1110111: c <= 9'b1001000;
				8'b101011: c <= 9'b11011;
				8'b1101011: c <= 9'b101101;
				8'b111100: c <= 9'b11101011;
				8'b1000111: c <= 9'b110110110;
				8'b1011111: c <= 9'b100000000;
				8'b1110100: c <= 9'b100101101;
				8'b101101: c <= 9'b1010111;
				8'b1010011: c <= 9'b100001100;
				8'b1100001: c <= 9'b10000;
				8'b110101: c <= 9'b1010110;
				8'b1000100: c <= 9'b110100000;
				8'b1010001: c <= 9'b11011110;
				8'b1010100: c <= 9'b101111001;
				8'b1100110: c <= 9'b111001010;
				8'b101010: c <= 9'b1110010;
				8'b1011110: c <= 9'b10101100;
				8'b1100111: c <= 9'b111000;
				8'b1011010: c <= 9'b111111010;
				8'b1000010: c <= 9'b110010001;
				8'b111101: c <= 9'b110101001;
				8'b110000: c <= 9'b110001101;
				8'b111110: c <= 9'b100011001;
				8'b1100010: c <= 9'b110000010;
				8'b1110000: c <= 9'b111011001;
				8'b1101001: c <= 9'b11110001;
				8'b1110011: c <= 9'b100101010;
				8'b1001100: c <= 9'b111100011;
				8'b100001: c <= 9'b11111101;
				8'b1000110: c <= 9'b11101000;
				8'b1110010: c <= 9'b1;
				8'b1010000: c <= 9'b11111011;
				8'b1111010: c <= 9'b1111100;
				8'b1010101: c <= 9'b110110010;
				8'b111011: c <= 9'b1000101;
				8'b1001101: c <= 9'b10000011;
				8'b111111: c <= 9'b11101000;
				8'b1101110: c <= 9'b1100000;
				8'b1111011: c <= 9'b111111111;
				8'b1001011: c <= 9'b111011011;
				8'b1101111: c <= 9'b111101010;
				8'b1101000: c <= 9'b11001010;
				8'b101100: c <= 9'b101001;
				8'b100100: c <= 9'b10110101;
				8'b1111000: c <= 9'b111111110;
				8'b1000101: c <= 9'b11100010;
				8'b1011001: c <= 9'b101100011;
				8'b110100: c <= 9'b11100010;
				8'b1111001: c <= 9'b110100100;
				8'b1110001: c <= 9'b100100000;
				8'b1001111: c <= 9'b10111111;
				8'b1100101: c <= 9'b10100100;
				8'b1111110: c <= 9'b111100001;
				8'b1111100: c <= 9'b110101011;
				8'b1010110: c <= 9'b110100000;
				8'b110010: c <= 9'b110100010;
				8'b1101101: c <= 9'b110111100;
				8'b100011: c <= 9'b101110011;
				8'b1110101: c <= 9'b1011000;
				8'b1111101: c <= 9'b100110011;
				8'b101001: c <= 9'b111000101;
				8'b1010010: c <= 9'b11110000;
				8'b1011000: c <= 9'b1001110;
				8'b101110: c <= 9'b111001101;
				8'b1000001: c <= 9'b10111101;
				default: c <= 9'b0;
			endcase
			9'b10110001 : case(di)
				8'b1000011: c <= 9'b110010011;
				8'b101000: c <= 9'b111000000;
				8'b111010: c <= 9'b10101011;
				8'b110110: c <= 9'b110010111;
				8'b1100100: c <= 9'b1111011;
				8'b1000000: c <= 9'b110101111;
				8'b1110110: c <= 9'b100111101;
				8'b100101: c <= 9'b110010100;
				8'b101111: c <= 9'b111110101;
				8'b100110: c <= 9'b110010010;
				8'b1100011: c <= 9'b100010101;
				8'b1001000: c <= 9'b100000111;
				8'b111000: c <= 9'b110000;
				8'b110001: c <= 9'b101101100;
				8'b1010111: c <= 9'b111011010;
				8'b1001110: c <= 9'b100010100;
				8'b1101010: c <= 9'b110111;
				8'b1001001: c <= 9'b100111101;
				8'b1100000: c <= 9'b11000111;
				8'b110111: c <= 9'b101000111;
				8'b1011101: c <= 9'b110000110;
				8'b1011011: c <= 9'b10110011;
				8'b111001: c <= 9'b110100011;
				8'b1001010: c <= 9'b111100111;
				8'b110011: c <= 9'b101010100;
				8'b1101100: c <= 9'b111011;
				8'b1110111: c <= 9'b1111000;
				8'b101011: c <= 9'b11110110;
				8'b1101011: c <= 9'b11010101;
				8'b111100: c <= 9'b110000011;
				8'b1000111: c <= 9'b10011010;
				8'b1011111: c <= 9'b111001011;
				8'b1110100: c <= 9'b101110010;
				8'b101101: c <= 9'b101000101;
				8'b1010011: c <= 9'b101110001;
				8'b1100001: c <= 9'b100011100;
				8'b110101: c <= 9'b111000011;
				8'b1000100: c <= 9'b111010111;
				8'b1010001: c <= 9'b110001001;
				8'b1010100: c <= 9'b101010000;
				8'b1100110: c <= 9'b100011101;
				8'b101010: c <= 9'b110000111;
				8'b1011110: c <= 9'b111101010;
				8'b1100111: c <= 9'b11111001;
				8'b1011010: c <= 9'b110110011;
				8'b1000010: c <= 9'b1001;
				8'b111101: c <= 9'b100110110;
				8'b110000: c <= 9'b110101111;
				8'b111110: c <= 9'b110100010;
				8'b1100010: c <= 9'b1100001;
				8'b1110000: c <= 9'b101000011;
				8'b1101001: c <= 9'b1001110;
				8'b1110011: c <= 9'b101111000;
				8'b1001100: c <= 9'b101111110;
				8'b100001: c <= 9'b111000111;
				8'b1000110: c <= 9'b111101110;
				8'b1110010: c <= 9'b1100000;
				8'b1010000: c <= 9'b10010111;
				8'b1111010: c <= 9'b101111000;
				8'b1010101: c <= 9'b10011000;
				8'b111011: c <= 9'b100000011;
				8'b1001101: c <= 9'b100110011;
				8'b111111: c <= 9'b100010011;
				8'b1101110: c <= 9'b101010111;
				8'b1111011: c <= 9'b110110100;
				8'b1001011: c <= 9'b1101110;
				8'b1101111: c <= 9'b1010010;
				8'b1101000: c <= 9'b100011000;
				8'b101100: c <= 9'b111000100;
				8'b100100: c <= 9'b1000101;
				8'b1111000: c <= 9'b101001010;
				8'b1000101: c <= 9'b11001111;
				8'b1011001: c <= 9'b110101;
				8'b110100: c <= 9'b10101010;
				8'b1111001: c <= 9'b111001010;
				8'b1110001: c <= 9'b101001010;
				8'b1001111: c <= 9'b100001101;
				8'b1100101: c <= 9'b1011111;
				8'b1111110: c <= 9'b110100110;
				8'b1111100: c <= 9'b11100010;
				8'b1010110: c <= 9'b11101;
				8'b110010: c <= 9'b100111101;
				8'b1101101: c <= 9'b111010111;
				8'b100011: c <= 9'b100001100;
				8'b1110101: c <= 9'b1010001;
				8'b1111101: c <= 9'b111001010;
				8'b101001: c <= 9'b110100100;
				8'b1010010: c <= 9'b101101111;
				8'b1011000: c <= 9'b10111011;
				8'b101110: c <= 9'b100101101;
				8'b1000001: c <= 9'b111010;
				default: c <= 9'b0;
			endcase
			9'b111101111 : case(di)
				8'b1000011: c <= 9'b100001110;
				8'b101000: c <= 9'b110110111;
				8'b111010: c <= 9'b100010100;
				8'b110110: c <= 9'b111100100;
				8'b1100100: c <= 9'b111101100;
				8'b1000000: c <= 9'b1100001;
				8'b1110110: c <= 9'b10111111;
				8'b100101: c <= 9'b101011010;
				8'b101111: c <= 9'b101110111;
				8'b100110: c <= 9'b101101110;
				8'b1100011: c <= 9'b1101100;
				8'b1001000: c <= 9'b111010000;
				8'b111000: c <= 9'b10010000;
				8'b110001: c <= 9'b111001;
				8'b1010111: c <= 9'b10011100;
				8'b1001110: c <= 9'b111010111;
				8'b1101010: c <= 9'b101;
				8'b1001001: c <= 9'b100011001;
				8'b1100000: c <= 9'b1111111;
				8'b110111: c <= 9'b101010101;
				8'b1011101: c <= 9'b11100100;
				8'b1011011: c <= 9'b10100110;
				8'b111001: c <= 9'b11011101;
				8'b1001010: c <= 9'b111010010;
				8'b110011: c <= 9'b11111100;
				8'b1101100: c <= 9'b100011111;
				8'b1110111: c <= 9'b101;
				8'b101011: c <= 9'b11100;
				8'b1101011: c <= 9'b100100000;
				8'b111100: c <= 9'b110001100;
				8'b1000111: c <= 9'b100100000;
				8'b1011111: c <= 9'b110111100;
				8'b1110100: c <= 9'b11101001;
				8'b101101: c <= 9'b100001100;
				8'b1010011: c <= 9'b11001;
				8'b1100001: c <= 9'b110011111;
				8'b110101: c <= 9'b101100000;
				8'b1000100: c <= 9'b111010010;
				8'b1010001: c <= 9'b110110010;
				8'b1010100: c <= 9'b1110010;
				8'b1100110: c <= 9'b100011100;
				8'b101010: c <= 9'b111011111;
				8'b1011110: c <= 9'b111000010;
				8'b1100111: c <= 9'b111000110;
				8'b1011010: c <= 9'b1111010;
				8'b1000010: c <= 9'b101101011;
				8'b111101: c <= 9'b1000011;
				8'b110000: c <= 9'b110011100;
				8'b111110: c <= 9'b110011001;
				8'b1100010: c <= 9'b100001010;
				8'b1110000: c <= 9'b1000100;
				8'b1101001: c <= 9'b10000110;
				8'b1110011: c <= 9'b10001011;
				8'b1001100: c <= 9'b110110;
				8'b100001: c <= 9'b1000;
				8'b1000110: c <= 9'b1100001;
				8'b1110010: c <= 9'b100110010;
				8'b1010000: c <= 9'b10101101;
				8'b1111010: c <= 9'b11000000;
				8'b1010101: c <= 9'b11001000;
				8'b111011: c <= 9'b100011;
				8'b1001101: c <= 9'b111;
				8'b111111: c <= 9'b11;
				8'b1101110: c <= 9'b111101000;
				8'b1111011: c <= 9'b111111010;
				8'b1001011: c <= 9'b110000010;
				8'b1101111: c <= 9'b10101100;
				8'b1101000: c <= 9'b111010111;
				8'b101100: c <= 9'b100010101;
				8'b100100: c <= 9'b111010010;
				8'b1111000: c <= 9'b1011111;
				8'b1000101: c <= 9'b11000011;
				8'b1011001: c <= 9'b10101100;
				8'b110100: c <= 9'b100110011;
				8'b1111001: c <= 9'b1010101;
				8'b1110001: c <= 9'b101011011;
				8'b1001111: c <= 9'b101010101;
				8'b1100101: c <= 9'b11100000;
				8'b1111110: c <= 9'b10011000;
				8'b1111100: c <= 9'b110111001;
				8'b1010110: c <= 9'b11010;
				8'b110010: c <= 9'b100110101;
				8'b1101101: c <= 9'b11101011;
				8'b100011: c <= 9'b10111111;
				8'b1110101: c <= 9'b101011001;
				8'b1111101: c <= 9'b11000000;
				8'b101001: c <= 9'b101011001;
				8'b1010010: c <= 9'b1111110;
				8'b1011000: c <= 9'b11110001;
				8'b101110: c <= 9'b111110001;
				8'b1000001: c <= 9'b1101101;
				default: c <= 9'b0;
			endcase
			9'b101110110 : case(di)
				8'b1000011: c <= 9'b1100001;
				8'b101000: c <= 9'b101100011;
				8'b111010: c <= 9'b110100101;
				8'b110110: c <= 9'b1001011;
				8'b1100100: c <= 9'b110011;
				8'b1000000: c <= 9'b10001011;
				8'b1110110: c <= 9'b11111011;
				8'b100101: c <= 9'b100;
				8'b101111: c <= 9'b1100100;
				8'b100110: c <= 9'b100100;
				8'b1100011: c <= 9'b101000110;
				8'b1001000: c <= 9'b111101111;
				8'b111000: c <= 9'b110010001;
				8'b110001: c <= 9'b101101001;
				8'b1010111: c <= 9'b10011001;
				8'b1001110: c <= 9'b100111101;
				8'b1101010: c <= 9'b1010110;
				8'b1001001: c <= 9'b10100;
				8'b1100000: c <= 9'b111101001;
				8'b110111: c <= 9'b11001011;
				8'b1011101: c <= 9'b100101101;
				8'b1011011: c <= 9'b11001;
				8'b111001: c <= 9'b11001000;
				8'b1001010: c <= 9'b101011110;
				8'b110011: c <= 9'b100010001;
				8'b1101100: c <= 9'b111100010;
				8'b1110111: c <= 9'b101111110;
				8'b101011: c <= 9'b11010010;
				8'b1101011: c <= 9'b11100;
				8'b111100: c <= 9'b101000001;
				8'b1000111: c <= 9'b101010100;
				8'b1011111: c <= 9'b101110110;
				8'b1110100: c <= 9'b11001010;
				8'b101101: c <= 9'b111000011;
				8'b1010011: c <= 9'b10000101;
				8'b1100001: c <= 9'b101011111;
				8'b110101: c <= 9'b10010000;
				8'b1000100: c <= 9'b10000010;
				8'b1010001: c <= 9'b11100110;
				8'b1010100: c <= 9'b10000011;
				8'b1100110: c <= 9'b11010000;
				8'b101010: c <= 9'b111;
				8'b1011110: c <= 9'b110101010;
				8'b1100111: c <= 9'b1100011;
				8'b1011010: c <= 9'b1101100;
				8'b1000010: c <= 9'b110000;
				8'b111101: c <= 9'b10000001;
				8'b110000: c <= 9'b1011011;
				8'b111110: c <= 9'b10011011;
				8'b1100010: c <= 9'b111111011;
				8'b1110000: c <= 9'b1011111;
				8'b1101001: c <= 9'b100101101;
				8'b1110011: c <= 9'b11110101;
				8'b1001100: c <= 9'b10000110;
				8'b100001: c <= 9'b1000110;
				8'b1000110: c <= 9'b1100010;
				8'b1110010: c <= 9'b110100000;
				8'b1010000: c <= 9'b11001010;
				8'b1111010: c <= 9'b1111001;
				8'b1010101: c <= 9'b1011000;
				8'b111011: c <= 9'b111011100;
				8'b1001101: c <= 9'b11100111;
				8'b111111: c <= 9'b101001;
				8'b1101110: c <= 9'b101100110;
				8'b1111011: c <= 9'b10010000;
				8'b1001011: c <= 9'b111100;
				8'b1101111: c <= 9'b101111010;
				8'b1101000: c <= 9'b100;
				8'b101100: c <= 9'b100111011;
				8'b100100: c <= 9'b11101001;
				8'b1111000: c <= 9'b10110010;
				8'b1000101: c <= 9'b110001;
				8'b1011001: c <= 9'b101000011;
				8'b110100: c <= 9'b101101110;
				8'b1111001: c <= 9'b100010110;
				8'b1110001: c <= 9'b101100000;
				8'b1001111: c <= 9'b1001100;
				8'b1100101: c <= 9'b1101101;
				8'b1111110: c <= 9'b10100000;
				8'b1111100: c <= 9'b111001001;
				8'b1010110: c <= 9'b10000001;
				8'b110010: c <= 9'b100011011;
				8'b1101101: c <= 9'b110100110;
				8'b100011: c <= 9'b111010010;
				8'b1110101: c <= 9'b11110110;
				8'b1111101: c <= 9'b11100110;
				8'b101001: c <= 9'b1011;
				8'b1010010: c <= 9'b100111001;
				8'b1011000: c <= 9'b101000100;
				8'b101110: c <= 9'b100000000;
				8'b1000001: c <= 9'b1100010;
				default: c <= 9'b0;
			endcase
			9'b101100110 : case(di)
				8'b1000011: c <= 9'b111100100;
				8'b101000: c <= 9'b110110100;
				8'b111010: c <= 9'b100011000;
				8'b110110: c <= 9'b100111;
				8'b1100100: c <= 9'b10100010;
				8'b1000000: c <= 9'b11011101;
				8'b1110110: c <= 9'b110001111;
				8'b100101: c <= 9'b10010000;
				8'b101111: c <= 9'b110000111;
				8'b100110: c <= 9'b101110111;
				8'b1100011: c <= 9'b1100111;
				8'b1001000: c <= 9'b100100111;
				8'b111000: c <= 9'b1001;
				8'b110001: c <= 9'b1011110;
				8'b1010111: c <= 9'b100011100;
				8'b1001110: c <= 9'b1000011;
				8'b1101010: c <= 9'b111101;
				8'b1001001: c <= 9'b110101011;
				8'b1100000: c <= 9'b110101101;
				8'b110111: c <= 9'b11100110;
				8'b1011101: c <= 9'b11101100;
				8'b1011011: c <= 9'b111011;
				8'b111001: c <= 9'b10010011;
				8'b1001010: c <= 9'b10000111;
				8'b110011: c <= 9'b100111011;
				8'b1101100: c <= 9'b1000;
				8'b1110111: c <= 9'b110001;
				8'b101011: c <= 9'b110010110;
				8'b1101011: c <= 9'b10101011;
				8'b111100: c <= 9'b110000001;
				8'b1000111: c <= 9'b11;
				8'b1011111: c <= 9'b110111010;
				8'b1110100: c <= 9'b110010001;
				8'b101101: c <= 9'b1111010;
				8'b1010011: c <= 9'b10001100;
				8'b1100001: c <= 9'b110000101;
				8'b110101: c <= 9'b10011;
				8'b1000100: c <= 9'b100101000;
				8'b1010001: c <= 9'b11000111;
				8'b1010100: c <= 9'b110110101;
				8'b1100110: c <= 9'b101010001;
				8'b101010: c <= 9'b100000010;
				8'b1011110: c <= 9'b11000111;
				8'b1100111: c <= 9'b111100101;
				8'b1011010: c <= 9'b11001101;
				8'b1000010: c <= 9'b101111010;
				8'b111101: c <= 9'b1110101;
				8'b110000: c <= 9'b111110011;
				8'b111110: c <= 9'b11100010;
				8'b1100010: c <= 9'b10010101;
				8'b1110000: c <= 9'b100111011;
				8'b1101001: c <= 9'b100101100;
				8'b1110011: c <= 9'b1011001;
				8'b1001100: c <= 9'b101100000;
				8'b100001: c <= 9'b111001101;
				8'b1000110: c <= 9'b10111100;
				8'b1110010: c <= 9'b111011001;
				8'b1010000: c <= 9'b1101100;
				8'b1111010: c <= 9'b1101101;
				8'b1010101: c <= 9'b101010011;
				8'b111011: c <= 9'b1111110;
				8'b1001101: c <= 9'b101100;
				8'b111111: c <= 9'b111011;
				8'b1101110: c <= 9'b1100110;
				8'b1111011: c <= 9'b11010101;
				8'b1001011: c <= 9'b11100001;
				8'b1101111: c <= 9'b101000011;
				8'b1101000: c <= 9'b101010100;
				8'b101100: c <= 9'b110000;
				8'b100100: c <= 9'b110001000;
				8'b1111000: c <= 9'b100110101;
				8'b1000101: c <= 9'b111000011;
				8'b1011001: c <= 9'b11100;
				8'b110100: c <= 9'b100101000;
				8'b1111001: c <= 9'b110110100;
				8'b1110001: c <= 9'b101;
				8'b1001111: c <= 9'b11001001;
				8'b1100101: c <= 9'b110001101;
				8'b1111110: c <= 9'b100000001;
				8'b1111100: c <= 9'b101111010;
				8'b1010110: c <= 9'b101110011;
				8'b110010: c <= 9'b10101111;
				8'b1101101: c <= 9'b110111;
				8'b100011: c <= 9'b11110111;
				8'b1110101: c <= 9'b10010110;
				8'b1111101: c <= 9'b100001010;
				8'b101001: c <= 9'b10110101;
				8'b1010010: c <= 9'b111010010;
				8'b1011000: c <= 9'b100101100;
				8'b101110: c <= 9'b11011011;
				8'b1000001: c <= 9'b111000110;
				default: c <= 9'b0;
			endcase
			9'b110011001 : case(di)
				8'b1000011: c <= 9'b110011111;
				8'b101000: c <= 9'b110011010;
				8'b111010: c <= 9'b101011111;
				8'b110110: c <= 9'b101011011;
				8'b1100100: c <= 9'b11111100;
				8'b1000000: c <= 9'b1111100;
				8'b1110110: c <= 9'b101001011;
				8'b100101: c <= 9'b10111011;
				8'b101111: c <= 9'b100100010;
				8'b100110: c <= 9'b111;
				8'b1100011: c <= 9'b111100110;
				8'b1001000: c <= 9'b100010110;
				8'b111000: c <= 9'b111001001;
				8'b110001: c <= 9'b100001010;
				8'b1010111: c <= 9'b10011001;
				8'b1001110: c <= 9'b100110;
				8'b1101010: c <= 9'b10001001;
				8'b1001001: c <= 9'b111010;
				8'b1100000: c <= 9'b111011010;
				8'b110111: c <= 9'b10011001;
				8'b1011101: c <= 9'b110101011;
				8'b1011011: c <= 9'b10010000;
				8'b111001: c <= 9'b1101101;
				8'b1001010: c <= 9'b11011001;
				8'b110011: c <= 9'b111001101;
				8'b1101100: c <= 9'b1011010;
				8'b1110111: c <= 9'b1110111;
				8'b101011: c <= 9'b11011010;
				8'b1101011: c <= 9'b111111010;
				8'b111100: c <= 9'b11111000;
				8'b1000111: c <= 9'b101000111;
				8'b1011111: c <= 9'b11000000;
				8'b1110100: c <= 9'b101011000;
				8'b101101: c <= 9'b111;
				8'b1010011: c <= 9'b1010001;
				8'b1100001: c <= 9'b10011001;
				8'b110101: c <= 9'b11100000;
				8'b1000100: c <= 9'b11000111;
				8'b1010001: c <= 9'b11100010;
				8'b1010100: c <= 9'b100001100;
				8'b1100110: c <= 9'b101001110;
				8'b101010: c <= 9'b100010110;
				8'b1011110: c <= 9'b100111100;
				8'b1100111: c <= 9'b1100101;
				8'b1011010: c <= 9'b11111000;
				8'b1000010: c <= 9'b11110011;
				8'b111101: c <= 9'b101010100;
				8'b110000: c <= 9'b100101011;
				8'b111110: c <= 9'b11001001;
				8'b1100010: c <= 9'b1111110;
				8'b1110000: c <= 9'b10101101;
				8'b1101001: c <= 9'b1101;
				8'b1110011: c <= 9'b101010;
				8'b1001100: c <= 9'b111111011;
				8'b100001: c <= 9'b100010000;
				8'b1000110: c <= 9'b10110111;
				8'b1110010: c <= 9'b100010011;
				8'b1010000: c <= 9'b1100100;
				8'b1111010: c <= 9'b11001110;
				8'b1010101: c <= 9'b110011110;
				8'b111011: c <= 9'b101100010;
				8'b1001101: c <= 9'b1010010;
				8'b111111: c <= 9'b10001001;
				8'b1101110: c <= 9'b110000011;
				8'b1111011: c <= 9'b110011110;
				8'b1001011: c <= 9'b101101100;
				8'b1101111: c <= 9'b110010001;
				8'b1101000: c <= 9'b100001010;
				8'b101100: c <= 9'b11110;
				8'b100100: c <= 9'b101001001;
				8'b1111000: c <= 9'b1001010;
				8'b1000101: c <= 9'b1000001;
				8'b1011001: c <= 9'b111111101;
				8'b110100: c <= 9'b100101000;
				8'b1111001: c <= 9'b101100011;
				8'b1110001: c <= 9'b100110101;
				8'b1001111: c <= 9'b110010;
				8'b1100101: c <= 9'b100001110;
				8'b1111110: c <= 9'b101000011;
				8'b1111100: c <= 9'b1100101;
				8'b1010110: c <= 9'b11100001;
				8'b110010: c <= 9'b100110111;
				8'b1101101: c <= 9'b111100011;
				8'b100011: c <= 9'b11010000;
				8'b1110101: c <= 9'b11101001;
				8'b1111101: c <= 9'b11100100;
				8'b101001: c <= 9'b11010011;
				8'b1010010: c <= 9'b10000101;
				8'b1011000: c <= 9'b111110001;
				8'b101110: c <= 9'b1011010;
				8'b1000001: c <= 9'b10000111;
				default: c <= 9'b0;
			endcase
			9'b100110 : case(di)
				8'b1000011: c <= 9'b10010110;
				8'b101000: c <= 9'b10000;
				8'b111010: c <= 9'b111001;
				8'b110110: c <= 9'b101001;
				8'b1100100: c <= 9'b11000000;
				8'b1000000: c <= 9'b101101011;
				8'b1110110: c <= 9'b1110010;
				8'b100101: c <= 9'b10110110;
				8'b101111: c <= 9'b110011110;
				8'b100110: c <= 9'b111000100;
				8'b1100011: c <= 9'b101101111;
				8'b1001000: c <= 9'b11011110;
				8'b111000: c <= 9'b110010010;
				8'b110001: c <= 9'b101000101;
				8'b1010111: c <= 9'b110111010;
				8'b1001110: c <= 9'b110010100;
				8'b1101010: c <= 9'b111110101;
				8'b1001001: c <= 9'b1111000;
				8'b1100000: c <= 9'b110110110;
				8'b110111: c <= 9'b11101111;
				8'b1011101: c <= 9'b1101111;
				8'b1011011: c <= 9'b11001010;
				8'b111001: c <= 9'b101110000;
				8'b1001010: c <= 9'b100011100;
				8'b110011: c <= 9'b10101010;
				8'b1101100: c <= 9'b101101000;
				8'b1110111: c <= 9'b10110;
				8'b101011: c <= 9'b110011011;
				8'b1101011: c <= 9'b110011010;
				8'b111100: c <= 9'b1100111;
				8'b1000111: c <= 9'b100000111;
				8'b1011111: c <= 9'b11001111;
				8'b1110100: c <= 9'b11101000;
				8'b101101: c <= 9'b11001101;
				8'b1010011: c <= 9'b110011010;
				8'b1100001: c <= 9'b11100001;
				8'b110101: c <= 9'b11110;
				8'b1000100: c <= 9'b100100101;
				8'b1010001: c <= 9'b11010;
				8'b1010100: c <= 9'b111110011;
				8'b1100110: c <= 9'b100101110;
				8'b101010: c <= 9'b100110100;
				8'b1011110: c <= 9'b10101101;
				8'b1100111: c <= 9'b110100010;
				8'b1011010: c <= 9'b100111111;
				8'b1000010: c <= 9'b111111000;
				8'b111101: c <= 9'b11110111;
				8'b110000: c <= 9'b10101110;
				8'b111110: c <= 9'b100100000;
				8'b1100010: c <= 9'b100110100;
				8'b1110000: c <= 9'b101110000;
				8'b1101001: c <= 9'b101011001;
				8'b1110011: c <= 9'b101110100;
				8'b1001100: c <= 9'b110000;
				8'b100001: c <= 9'b110001111;
				8'b1000110: c <= 9'b111100011;
				8'b1110010: c <= 9'b110011101;
				8'b1010000: c <= 9'b100101;
				8'b1111010: c <= 9'b1110001;
				8'b1010101: c <= 9'b100010111;
				8'b111011: c <= 9'b101101101;
				8'b1001101: c <= 9'b100011000;
				8'b111111: c <= 9'b101011011;
				8'b1101110: c <= 9'b100011000;
				8'b1111011: c <= 9'b111001101;
				8'b1001011: c <= 9'b111011110;
				8'b1101111: c <= 9'b10000010;
				8'b1101000: c <= 9'b100000010;
				8'b101100: c <= 9'b1000100;
				8'b100100: c <= 9'b101001;
				8'b1111000: c <= 9'b111110000;
				8'b1000101: c <= 9'b10100100;
				8'b1011001: c <= 9'b100010010;
				8'b110100: c <= 9'b10100110;
				8'b1111001: c <= 9'b110011011;
				8'b1110001: c <= 9'b11000111;
				8'b1001111: c <= 9'b1100110;
				8'b1100101: c <= 9'b100010111;
				8'b1111110: c <= 9'b111101101;
				8'b1111100: c <= 9'b100101010;
				8'b1010110: c <= 9'b11001;
				8'b110010: c <= 9'b101110011;
				8'b1101101: c <= 9'b11110110;
				8'b100011: c <= 9'b110000001;
				8'b1110101: c <= 9'b111101010;
				8'b1111101: c <= 9'b100101011;
				8'b101001: c <= 9'b10001110;
				8'b1010010: c <= 9'b100111111;
				8'b1011000: c <= 9'b111001010;
				8'b101110: c <= 9'b101101000;
				8'b1000001: c <= 9'b1000011;
				default: c <= 9'b0;
			endcase
			9'b110010100 : case(di)
				8'b1000011: c <= 9'b101110000;
				8'b101000: c <= 9'b101101101;
				8'b111010: c <= 9'b11110011;
				8'b110110: c <= 9'b111011001;
				8'b1100100: c <= 9'b1111011;
				8'b1000000: c <= 9'b1010111;
				8'b1110110: c <= 9'b101110001;
				8'b100101: c <= 9'b10100101;
				8'b101111: c <= 9'b100100010;
				8'b100110: c <= 9'b10100100;
				8'b1100011: c <= 9'b110011011;
				8'b1001000: c <= 9'b11011;
				8'b111000: c <= 9'b100011101;
				8'b110001: c <= 9'b100101000;
				8'b1010111: c <= 9'b10001110;
				8'b1001110: c <= 9'b1100011;
				8'b1101010: c <= 9'b100000100;
				8'b1001001: c <= 9'b10101111;
				8'b1100000: c <= 9'b1101001;
				8'b110111: c <= 9'b100111;
				8'b1011101: c <= 9'b100111101;
				8'b1011011: c <= 9'b11110010;
				8'b111001: c <= 9'b1111001;
				8'b1001010: c <= 9'b11111110;
				8'b110011: c <= 9'b110000101;
				8'b1101100: c <= 9'b1110011;
				8'b1110111: c <= 9'b111001001;
				8'b101011: c <= 9'b1010000;
				8'b1101011: c <= 9'b1100110;
				8'b111100: c <= 9'b101000011;
				8'b1000111: c <= 9'b10001001;
				8'b1011111: c <= 9'b1111;
				8'b1110100: c <= 9'b111101110;
				8'b101101: c <= 9'b100001011;
				8'b1010011: c <= 9'b110000110;
				8'b1100001: c <= 9'b111000110;
				8'b110101: c <= 9'b1001100;
				8'b1000100: c <= 9'b100;
				8'b1010001: c <= 9'b101000001;
				8'b1010100: c <= 9'b101110001;
				8'b1100110: c <= 9'b11010010;
				8'b101010: c <= 9'b11010001;
				8'b1011110: c <= 9'b10001001;
				8'b1100111: c <= 9'b101110100;
				8'b1011010: c <= 9'b111000100;
				8'b1000010: c <= 9'b10000110;
				8'b111101: c <= 9'b101110001;
				8'b110000: c <= 9'b100010;
				8'b111110: c <= 9'b10101000;
				8'b1100010: c <= 9'b101011110;
				8'b1110000: c <= 9'b100100110;
				8'b1101001: c <= 9'b101001110;
				8'b1110011: c <= 9'b1110000;
				8'b1001100: c <= 9'b111001111;
				8'b100001: c <= 9'b101000011;
				8'b1000110: c <= 9'b110011011;
				8'b1110010: c <= 9'b110110010;
				8'b1010000: c <= 9'b111000010;
				8'b1111010: c <= 9'b111010000;
				8'b1010101: c <= 9'b111111000;
				8'b111011: c <= 9'b100010010;
				8'b1001101: c <= 9'b110101011;
				8'b111111: c <= 9'b110111;
				8'b1101110: c <= 9'b101110010;
				8'b1111011: c <= 9'b11100000;
				8'b1001011: c <= 9'b100110111;
				8'b1101111: c <= 9'b110101;
				8'b1101000: c <= 9'b101110001;
				8'b101100: c <= 9'b111011110;
				8'b100100: c <= 9'b100100110;
				8'b1111000: c <= 9'b111100101;
				8'b1000101: c <= 9'b1111001;
				8'b1011001: c <= 9'b11001011;
				8'b110100: c <= 9'b101011000;
				8'b1111001: c <= 9'b101001000;
				8'b1110001: c <= 9'b101010111;
				8'b1001111: c <= 9'b110101101;
				8'b1100101: c <= 9'b110000101;
				8'b1111110: c <= 9'b1010010;
				8'b1111100: c <= 9'b101101011;
				8'b1010110: c <= 9'b111011010;
				8'b110010: c <= 9'b110110111;
				8'b1101101: c <= 9'b1000110;
				8'b100011: c <= 9'b101010111;
				8'b1110101: c <= 9'b101011001;
				8'b1111101: c <= 9'b110110011;
				8'b101001: c <= 9'b110000000;
				8'b1010010: c <= 9'b110101011;
				8'b1011000: c <= 9'b111101100;
				8'b101110: c <= 9'b101110101;
				8'b1000001: c <= 9'b100011001;
				default: c <= 9'b0;
			endcase
			9'b110100100 : case(di)
				8'b1000011: c <= 9'b11100101;
				8'b101000: c <= 9'b10110011;
				8'b111010: c <= 9'b1110111;
				8'b110110: c <= 9'b101101010;
				8'b1100100: c <= 9'b10001010;
				8'b1000000: c <= 9'b11000000;
				8'b1110110: c <= 9'b110111100;
				8'b100101: c <= 9'b101011010;
				8'b101111: c <= 9'b1000110;
				8'b100110: c <= 9'b110011;
				8'b1100011: c <= 9'b111001101;
				8'b1001000: c <= 9'b1010010;
				8'b111000: c <= 9'b1011000;
				8'b110001: c <= 9'b111001010;
				8'b1010111: c <= 9'b1110000;
				8'b1001110: c <= 9'b1001100;
				8'b1101010: c <= 9'b1100001;
				8'b1001001: c <= 9'b11110100;
				8'b1100000: c <= 9'b11010111;
				8'b110111: c <= 9'b1010110;
				8'b1011101: c <= 9'b100111111;
				8'b1011011: c <= 9'b10010;
				8'b111001: c <= 9'b1011000;
				8'b1001010: c <= 9'b11110111;
				8'b110011: c <= 9'b101101001;
				8'b1101100: c <= 9'b110111;
				8'b1110111: c <= 9'b10110010;
				8'b101011: c <= 9'b101010010;
				8'b1101011: c <= 9'b100111010;
				8'b111100: c <= 9'b100101000;
				8'b1000111: c <= 9'b1000;
				8'b1011111: c <= 9'b11001000;
				8'b1110100: c <= 9'b11110100;
				8'b101101: c <= 9'b10000011;
				8'b1010011: c <= 9'b100000001;
				8'b1100001: c <= 9'b11;
				8'b110101: c <= 9'b111101001;
				8'b1000100: c <= 9'b10;
				8'b1010001: c <= 9'b11000100;
				8'b1010100: c <= 9'b10111011;
				8'b1100110: c <= 9'b101000101;
				8'b101010: c <= 9'b1001000;
				8'b1011110: c <= 9'b10011000;
				8'b1100111: c <= 9'b110100010;
				8'b1011010: c <= 9'b110000101;
				8'b1000010: c <= 9'b111011;
				8'b111101: c <= 9'b100010111;
				8'b110000: c <= 9'b101001010;
				8'b111110: c <= 9'b100001001;
				8'b1100010: c <= 9'b11111000;
				8'b1110000: c <= 9'b100001111;
				8'b1101001: c <= 9'b10111000;
				8'b1110011: c <= 9'b100101111;
				8'b1001100: c <= 9'b110100000;
				8'b100001: c <= 9'b101000111;
				8'b1000110: c <= 9'b10111111;
				8'b1110010: c <= 9'b10011;
				8'b1010000: c <= 9'b11010111;
				8'b1111010: c <= 9'b111011100;
				8'b1010101: c <= 9'b1010111;
				8'b111011: c <= 9'b1100;
				8'b1001101: c <= 9'b110000;
				8'b111111: c <= 9'b10101100;
				8'b1101110: c <= 9'b101101101;
				8'b1111011: c <= 9'b1010110;
				8'b1001011: c <= 9'b101011110;
				8'b1101111: c <= 9'b101100010;
				8'b1101000: c <= 9'b10100101;
				8'b101100: c <= 9'b10000010;
				8'b100100: c <= 9'b100001101;
				8'b1111000: c <= 9'b100110111;
				8'b1000101: c <= 9'b101000100;
				8'b1011001: c <= 9'b101011000;
				8'b110100: c <= 9'b101011110;
				8'b1111001: c <= 9'b100110010;
				8'b1110001: c <= 9'b111100110;
				8'b1001111: c <= 9'b1100100;
				8'b1100101: c <= 9'b110000010;
				8'b1111110: c <= 9'b101;
				8'b1111100: c <= 9'b101101000;
				8'b1010110: c <= 9'b101110010;
				8'b110010: c <= 9'b100011101;
				8'b1101101: c <= 9'b10110;
				8'b100011: c <= 9'b110000010;
				8'b1110101: c <= 9'b10110101;
				8'b1111101: c <= 9'b101000;
				8'b101001: c <= 9'b100001100;
				8'b1010010: c <= 9'b100111110;
				8'b1011000: c <= 9'b100010111;
				8'b101110: c <= 9'b10001110;
				8'b1000001: c <= 9'b11011;
				default: c <= 9'b0;
			endcase
			9'b1000000 : case(di)
				8'b1000011: c <= 9'b110000000;
				8'b101000: c <= 9'b101110001;
				8'b111010: c <= 9'b100000101;
				8'b110110: c <= 9'b110001000;
				8'b1100100: c <= 9'b1001011;
				8'b1000000: c <= 9'b11100111;
				8'b1110110: c <= 9'b110110;
				8'b100101: c <= 9'b100100;
				8'b101111: c <= 9'b101110;
				8'b100110: c <= 9'b101011000;
				8'b1100011: c <= 9'b101011;
				8'b1001000: c <= 9'b11001110;
				8'b111000: c <= 9'b110110000;
				8'b110001: c <= 9'b110010111;
				8'b1010111: c <= 9'b1001011;
				8'b1001110: c <= 9'b101001010;
				8'b1101010: c <= 9'b100110100;
				8'b1001001: c <= 9'b101101111;
				8'b1100000: c <= 9'b101000;
				8'b110111: c <= 9'b110101001;
				8'b1011101: c <= 9'b111110110;
				8'b1011011: c <= 9'b11110110;
				8'b111001: c <= 9'b100011000;
				8'b1001010: c <= 9'b10110111;
				8'b110011: c <= 9'b10001011;
				8'b1101100: c <= 9'b1100101;
				8'b1110111: c <= 9'b101010011;
				8'b101011: c <= 9'b111010110;
				8'b1101011: c <= 9'b110011000;
				8'b111100: c <= 9'b101111111;
				8'b1000111: c <= 9'b100111110;
				8'b1011111: c <= 9'b10110011;
				8'b1110100: c <= 9'b11100101;
				8'b101101: c <= 9'b100100011;
				8'b1010011: c <= 9'b11100000;
				8'b1100001: c <= 9'b10101101;
				8'b110101: c <= 9'b1111010;
				8'b1000100: c <= 9'b101001001;
				8'b1010001: c <= 9'b10001111;
				8'b1010100: c <= 9'b110011100;
				8'b1100110: c <= 9'b11010010;
				8'b101010: c <= 9'b11111101;
				8'b1011110: c <= 9'b10101000;
				8'b1100111: c <= 9'b100100010;
				8'b1011010: c <= 9'b11000011;
				8'b1000010: c <= 9'b101101100;
				8'b111101: c <= 9'b110001011;
				8'b110000: c <= 9'b11100101;
				8'b111110: c <= 9'b110011001;
				8'b1100010: c <= 9'b100111010;
				8'b1110000: c <= 9'b11111001;
				8'b1101001: c <= 9'b100001100;
				8'b1110011: c <= 9'b110000010;
				8'b1001100: c <= 9'b111100011;
				8'b100001: c <= 9'b10110101;
				8'b1000110: c <= 9'b110100011;
				8'b1110010: c <= 9'b111011101;
				8'b1010000: c <= 9'b11110111;
				8'b1111010: c <= 9'b111010010;
				8'b1010101: c <= 9'b10111;
				8'b111011: c <= 9'b11100011;
				8'b1001101: c <= 9'b1001110;
				8'b111111: c <= 9'b10100000;
				8'b1101110: c <= 9'b100110100;
				8'b1111011: c <= 9'b111110000;
				8'b1001011: c <= 9'b11011;
				8'b1101111: c <= 9'b111101000;
				8'b1101000: c <= 9'b100010010;
				8'b101100: c <= 9'b111111101;
				8'b100100: c <= 9'b100001110;
				8'b1111000: c <= 9'b1110100;
				8'b1000101: c <= 9'b11111000;
				8'b1011001: c <= 9'b110101010;
				8'b110100: c <= 9'b10110011;
				8'b1111001: c <= 9'b11001111;
				8'b1110001: c <= 9'b11000100;
				8'b1001111: c <= 9'b110110;
				8'b1100101: c <= 9'b111000100;
				8'b1111110: c <= 9'b111101010;
				8'b1111100: c <= 9'b111011010;
				8'b1010110: c <= 9'b110101010;
				8'b110010: c <= 9'b101111111;
				8'b1101101: c <= 9'b11000000;
				8'b100011: c <= 9'b1011111;
				8'b1110101: c <= 9'b10111010;
				8'b1111101: c <= 9'b1000010;
				8'b101001: c <= 9'b100010;
				8'b1010010: c <= 9'b101010011;
				8'b1011000: c <= 9'b11101000;
				8'b101110: c <= 9'b10011010;
				8'b1000001: c <= 9'b11110111;
				default: c <= 9'b0;
			endcase
			9'b1011 : case(di)
				8'b1000011: c <= 9'b1111000;
				8'b101000: c <= 9'b110100000;
				8'b111010: c <= 9'b101100;
				8'b110110: c <= 9'b10111011;
				8'b1100100: c <= 9'b11101111;
				8'b1000000: c <= 9'b110100001;
				8'b1110110: c <= 9'b10101001;
				8'b100101: c <= 9'b10011011;
				8'b101111: c <= 9'b110111110;
				8'b100110: c <= 9'b1000100;
				8'b1100011: c <= 9'b10001101;
				8'b1001000: c <= 9'b11000100;
				8'b111000: c <= 9'b101010100;
				8'b110001: c <= 9'b111110000;
				8'b1010111: c <= 9'b101101111;
				8'b1001110: c <= 9'b100101101;
				8'b1101010: c <= 9'b10110001;
				8'b1001001: c <= 9'b1000010;
				8'b1100000: c <= 9'b1010000;
				8'b110111: c <= 9'b110000110;
				8'b1011101: c <= 9'b11110101;
				8'b1011011: c <= 9'b101110000;
				8'b111001: c <= 9'b1110000;
				8'b1001010: c <= 9'b11000001;
				8'b110011: c <= 9'b100110100;
				8'b1101100: c <= 9'b10101110;
				8'b1110111: c <= 9'b110101010;
				8'b101011: c <= 9'b1010101;
				8'b1101011: c <= 9'b100010101;
				8'b111100: c <= 9'b110110100;
				8'b1000111: c <= 9'b1100100;
				8'b1011111: c <= 9'b1101111;
				8'b1110100: c <= 9'b111010111;
				8'b101101: c <= 9'b10000010;
				8'b1010011: c <= 9'b1010111;
				8'b1100001: c <= 9'b1001110;
				8'b110101: c <= 9'b110011011;
				8'b1000100: c <= 9'b110110010;
				8'b1010001: c <= 9'b110001011;
				8'b1010100: c <= 9'b11110101;
				8'b1100110: c <= 9'b111011100;
				8'b101010: c <= 9'b110110011;
				8'b1011110: c <= 9'b101010011;
				8'b1100111: c <= 9'b1000110;
				8'b1011010: c <= 9'b1110101;
				8'b1000010: c <= 9'b11011101;
				8'b111101: c <= 9'b110011000;
				8'b110000: c <= 9'b10000000;
				8'b111110: c <= 9'b1011100;
				8'b1100010: c <= 9'b110010001;
				8'b1110000: c <= 9'b11011100;
				8'b1101001: c <= 9'b1101100;
				8'b1110011: c <= 9'b11100000;
				8'b1001100: c <= 9'b11111100;
				8'b100001: c <= 9'b10011011;
				8'b1000110: c <= 9'b101101;
				8'b1110010: c <= 9'b101101110;
				8'b1010000: c <= 9'b10010101;
				8'b1111010: c <= 9'b10011011;
				8'b1010101: c <= 9'b1101010;
				8'b111011: c <= 9'b1101010;
				8'b1001101: c <= 9'b100111001;
				8'b111111: c <= 9'b101111000;
				8'b1101110: c <= 9'b11000011;
				8'b1111011: c <= 9'b110100010;
				8'b1001011: c <= 9'b111001111;
				8'b1101111: c <= 9'b1011111;
				8'b1101000: c <= 9'b10100010;
				8'b101100: c <= 9'b111100001;
				8'b100100: c <= 9'b111011010;
				8'b1111000: c <= 9'b111001101;
				8'b1000101: c <= 9'b11011000;
				8'b1011001: c <= 9'b110010011;
				8'b110100: c <= 9'b101011011;
				8'b1111001: c <= 9'b101011000;
				8'b1110001: c <= 9'b111101000;
				8'b1001111: c <= 9'b1001110;
				8'b1100101: c <= 9'b11000010;
				8'b1111110: c <= 9'b101110110;
				8'b1111100: c <= 9'b11101001;
				8'b1010110: c <= 9'b100001110;
				8'b110010: c <= 9'b100001111;
				8'b1101101: c <= 9'b101011101;
				8'b100011: c <= 9'b100110;
				8'b1110101: c <= 9'b111101101;
				8'b1111101: c <= 9'b100101101;
				8'b101001: c <= 9'b1110010;
				8'b1010010: c <= 9'b10100;
				8'b1011000: c <= 9'b10011100;
				8'b101110: c <= 9'b1010000;
				8'b1000001: c <= 9'b11001110;
				default: c <= 9'b0;
			endcase
			9'b1001100 : case(di)
				8'b1000011: c <= 9'b110101010;
				8'b101000: c <= 9'b111010000;
				8'b111010: c <= 9'b111010111;
				8'b110110: c <= 9'b110100001;
				8'b1100100: c <= 9'b1100000;
				8'b1000000: c <= 9'b11001000;
				8'b1110110: c <= 9'b11110;
				8'b100101: c <= 9'b11110110;
				8'b101111: c <= 9'b111111101;
				8'b100110: c <= 9'b100001;
				8'b1100011: c <= 9'b110001011;
				8'b1001000: c <= 9'b101110111;
				8'b111000: c <= 9'b111111000;
				8'b110001: c <= 9'b100101;
				8'b1010111: c <= 9'b1110000;
				8'b1001110: c <= 9'b111111101;
				8'b1101010: c <= 9'b100111001;
				8'b1001001: c <= 9'b101000101;
				8'b1100000: c <= 9'b1111001;
				8'b110111: c <= 9'b11111011;
				8'b1011101: c <= 9'b10001100;
				8'b1011011: c <= 9'b110101100;
				8'b111001: c <= 9'b100001011;
				8'b1001010: c <= 9'b1101100;
				8'b110011: c <= 9'b110011101;
				8'b1101100: c <= 9'b1101010;
				8'b1110111: c <= 9'b111011101;
				8'b101011: c <= 9'b111001100;
				8'b1101011: c <= 9'b110111110;
				8'b111100: c <= 9'b11111011;
				8'b1000111: c <= 9'b11000010;
				8'b1011111: c <= 9'b10010;
				8'b1110100: c <= 9'b100101000;
				8'b101101: c <= 9'b10001001;
				8'b1010011: c <= 9'b111101010;
				8'b1100001: c <= 9'b111011010;
				8'b110101: c <= 9'b10111001;
				8'b1000100: c <= 9'b10011;
				8'b1010001: c <= 9'b111110011;
				8'b1010100: c <= 9'b1011111;
				8'b1100110: c <= 9'b11000100;
				8'b101010: c <= 9'b11011110;
				8'b1011110: c <= 9'b110111011;
				8'b1100111: c <= 9'b1100110;
				8'b1011010: c <= 9'b1100101;
				8'b1000010: c <= 9'b1000100;
				8'b111101: c <= 9'b100101010;
				8'b110000: c <= 9'b11000010;
				8'b111110: c <= 9'b1101100;
				8'b1100010: c <= 9'b10101011;
				8'b1110000: c <= 9'b110000;
				8'b1101001: c <= 9'b1111101;
				8'b1110011: c <= 9'b110011000;
				8'b1001100: c <= 9'b101000101;
				8'b100001: c <= 9'b1110011;
				8'b1000110: c <= 9'b11100100;
				8'b1110010: c <= 9'b1011;
				8'b1010000: c <= 9'b11101111;
				8'b1111010: c <= 9'b111001001;
				8'b1010101: c <= 9'b111;
				8'b111011: c <= 9'b101011000;
				8'b1001101: c <= 9'b100101110;
				8'b111111: c <= 9'b10101111;
				8'b1101110: c <= 9'b10101110;
				8'b1111011: c <= 9'b110100110;
				8'b1001011: c <= 9'b101111001;
				8'b1101111: c <= 9'b101001011;
				8'b1101000: c <= 9'b110011010;
				8'b101100: c <= 9'b101110110;
				8'b100100: c <= 9'b110110111;
				8'b1111000: c <= 9'b1100010;
				8'b1000101: c <= 9'b101100110;
				8'b1011001: c <= 9'b110010101;
				8'b110100: c <= 9'b110010010;
				8'b1111001: c <= 9'b11010100;
				8'b1110001: c <= 9'b110001111;
				8'b1001111: c <= 9'b10001000;
				8'b1100101: c <= 9'b11100011;
				8'b1111110: c <= 9'b110111;
				8'b1111100: c <= 9'b101011000;
				8'b1010110: c <= 9'b10111001;
				8'b110010: c <= 9'b111111110;
				8'b1101101: c <= 9'b10011100;
				8'b100011: c <= 9'b110010011;
				8'b1110101: c <= 9'b101011000;
				8'b1111101: c <= 9'b111001001;
				8'b101001: c <= 9'b111110011;
				8'b1010010: c <= 9'b10111011;
				8'b1011000: c <= 9'b11010011;
				8'b101110: c <= 9'b11100111;
				8'b1000001: c <= 9'b110000011;
				default: c <= 9'b0;
			endcase
			9'b10010001 : case(di)
				8'b1000011: c <= 9'b101100100;
				8'b101000: c <= 9'b110010101;
				8'b111010: c <= 9'b11110111;
				8'b110110: c <= 9'b1101010;
				8'b1100100: c <= 9'b1000110;
				8'b1000000: c <= 9'b111001110;
				8'b1110110: c <= 9'b1001000;
				8'b100101: c <= 9'b101010100;
				8'b101111: c <= 9'b100000110;
				8'b100110: c <= 9'b101010010;
				8'b1100011: c <= 9'b11111;
				8'b1001000: c <= 9'b100101011;
				8'b111000: c <= 9'b10111011;
				8'b110001: c <= 9'b111011010;
				8'b1010111: c <= 9'b10010101;
				8'b1001110: c <= 9'b101110000;
				8'b1101010: c <= 9'b1000000;
				8'b1001001: c <= 9'b11010000;
				8'b1100000: c <= 9'b110011111;
				8'b110111: c <= 9'b11100100;
				8'b1011101: c <= 9'b11110100;
				8'b1011011: c <= 9'b100000101;
				8'b111001: c <= 9'b11101111;
				8'b1001010: c <= 9'b11001001;
				8'b110011: c <= 9'b10100111;
				8'b1101100: c <= 9'b100100110;
				8'b1110111: c <= 9'b1000001;
				8'b101011: c <= 9'b100101010;
				8'b1101011: c <= 9'b100001011;
				8'b111100: c <= 9'b11101;
				8'b1000111: c <= 9'b11100001;
				8'b1011111: c <= 9'b111001101;
				8'b1110100: c <= 9'b110110011;
				8'b101101: c <= 9'b110001;
				8'b1010011: c <= 9'b101011011;
				8'b1100001: c <= 9'b110011110;
				8'b110101: c <= 9'b100001100;
				8'b1000100: c <= 9'b100001001;
				8'b1010001: c <= 9'b1011011;
				8'b1010100: c <= 9'b101110001;
				8'b1100110: c <= 9'b10111011;
				8'b101010: c <= 9'b11011101;
				8'b1011110: c <= 9'b110110011;
				8'b1100111: c <= 9'b111100010;
				8'b1011010: c <= 9'b10000011;
				8'b1000010: c <= 9'b101001001;
				8'b111101: c <= 9'b111010000;
				8'b110000: c <= 9'b111001100;
				8'b111110: c <= 9'b11001111;
				8'b1100010: c <= 9'b100111;
				8'b1110000: c <= 9'b10010000;
				8'b1101001: c <= 9'b10111000;
				8'b1110011: c <= 9'b11111110;
				8'b1001100: c <= 9'b101001000;
				8'b100001: c <= 9'b11001001;
				8'b1000110: c <= 9'b111010000;
				8'b1110010: c <= 9'b1101110;
				8'b1010000: c <= 9'b111010001;
				8'b1111010: c <= 9'b10010001;
				8'b1010101: c <= 9'b100110;
				8'b111011: c <= 9'b100101101;
				8'b1001101: c <= 9'b101;
				8'b111111: c <= 9'b10001111;
				8'b1101110: c <= 9'b100000101;
				8'b1111011: c <= 9'b110011011;
				8'b1001011: c <= 9'b111111010;
				8'b1101111: c <= 9'b111101;
				8'b1101000: c <= 9'b100101001;
				8'b101100: c <= 9'b110001110;
				8'b100100: c <= 9'b11001110;
				8'b1111000: c <= 9'b1010011;
				8'b1000101: c <= 9'b110000111;
				8'b1011001: c <= 9'b11001011;
				8'b110100: c <= 9'b110010001;
				8'b1111001: c <= 9'b1101001;
				8'b1110001: c <= 9'b1000101;
				8'b1001111: c <= 9'b11110111;
				8'b1100101: c <= 9'b1111010;
				8'b1111110: c <= 9'b110111000;
				8'b1111100: c <= 9'b111101;
				8'b1010110: c <= 9'b11111;
				8'b110010: c <= 9'b101001111;
				8'b1101101: c <= 9'b10100101;
				8'b100011: c <= 9'b110001001;
				8'b1110101: c <= 9'b10011001;
				8'b1111101: c <= 9'b111101100;
				8'b101001: c <= 9'b10111000;
				8'b1010010: c <= 9'b100010011;
				8'b1011000: c <= 9'b100010011;
				8'b101110: c <= 9'b110001010;
				8'b1000001: c <= 9'b1110101;
				default: c <= 9'b0;
			endcase
			9'b100010001 : case(di)
				8'b1000011: c <= 9'b1110101;
				8'b101000: c <= 9'b101111111;
				8'b111010: c <= 9'b110101001;
				8'b110110: c <= 9'b11101000;
				8'b1100100: c <= 9'b10101001;
				8'b1000000: c <= 9'b10001100;
				8'b1110110: c <= 9'b111011100;
				8'b100101: c <= 9'b110010010;
				8'b101111: c <= 9'b101100010;
				8'b100110: c <= 9'b100000001;
				8'b1100011: c <= 9'b10001001;
				8'b1001000: c <= 9'b1100011;
				8'b111000: c <= 9'b101001011;
				8'b110001: c <= 9'b110111111;
				8'b1010111: c <= 9'b111000010;
				8'b1001110: c <= 9'b100110110;
				8'b1101010: c <= 9'b101100;
				8'b1001001: c <= 9'b100000110;
				8'b1100000: c <= 9'b110100000;
				8'b110111: c <= 9'b100010011;
				8'b1011101: c <= 9'b100111010;
				8'b1011011: c <= 9'b1001010;
				8'b111001: c <= 9'b100100110;
				8'b1001010: c <= 9'b1011111;
				8'b110011: c <= 9'b1010000;
				8'b1101100: c <= 9'b101100010;
				8'b1110111: c <= 9'b1110011;
				8'b101011: c <= 9'b1010010;
				8'b1101011: c <= 9'b11010100;
				8'b111100: c <= 9'b101011111;
				8'b1000111: c <= 9'b1000100;
				8'b1011111: c <= 9'b10111010;
				8'b1110100: c <= 9'b11110110;
				8'b101101: c <= 9'b11101111;
				8'b1010011: c <= 9'b11100110;
				8'b1100001: c <= 9'b10000001;
				8'b110101: c <= 9'b111000110;
				8'b1000100: c <= 9'b110000111;
				8'b1010001: c <= 9'b100100110;
				8'b1010100: c <= 9'b11110101;
				8'b1100110: c <= 9'b110011000;
				8'b101010: c <= 9'b11110000;
				8'b1011110: c <= 9'b10001011;
				8'b1100111: c <= 9'b111100101;
				8'b1011010: c <= 9'b11101111;
				8'b1000010: c <= 9'b100001110;
				8'b111101: c <= 9'b101000110;
				8'b110000: c <= 9'b1100100;
				8'b111110: c <= 9'b110100;
				8'b1100010: c <= 9'b110011100;
				8'b1110000: c <= 9'b11101011;
				8'b1101001: c <= 9'b11000110;
				8'b1110011: c <= 9'b11010011;
				8'b1001100: c <= 9'b11001011;
				8'b100001: c <= 9'b101000001;
				8'b1000110: c <= 9'b100001;
				8'b1110010: c <= 9'b100001100;
				8'b1010000: c <= 9'b1110;
				8'b1111010: c <= 9'b111111010;
				8'b1010101: c <= 9'b110001101;
				8'b111011: c <= 9'b110100010;
				8'b1001101: c <= 9'b111111110;
				8'b111111: c <= 9'b10011011;
				8'b1101110: c <= 9'b110001010;
				8'b1111011: c <= 9'b111111110;
				8'b1001011: c <= 9'b110011001;
				8'b1101111: c <= 9'b101;
				8'b1101000: c <= 9'b101101;
				8'b101100: c <= 9'b100011000;
				8'b100100: c <= 9'b110011000;
				8'b1111000: c <= 9'b101001110;
				8'b1000101: c <= 9'b11101111;
				8'b1011001: c <= 9'b110010100;
				8'b110100: c <= 9'b110111;
				8'b1111001: c <= 9'b10101000;
				8'b1110001: c <= 9'b11110110;
				8'b1001111: c <= 9'b1111101;
				8'b1100101: c <= 9'b111100111;
				8'b1111110: c <= 9'b101010100;
				8'b1111100: c <= 9'b110010101;
				8'b1010110: c <= 9'b10000111;
				8'b110010: c <= 9'b1111101;
				8'b1101101: c <= 9'b1000011;
				8'b100011: c <= 9'b111110110;
				8'b1110101: c <= 9'b110011001;
				8'b1111101: c <= 9'b110010010;
				8'b101001: c <= 9'b100100110;
				8'b1010010: c <= 9'b10011011;
				8'b1011000: c <= 9'b100001110;
				8'b101110: c <= 9'b110101001;
				8'b1000001: c <= 9'b10010111;
				default: c <= 9'b0;
			endcase
			9'b110100111 : case(di)
				8'b1000011: c <= 9'b101;
				8'b101000: c <= 9'b110110111;
				8'b111010: c <= 9'b10111011;
				8'b110110: c <= 9'b110001001;
				8'b1100100: c <= 9'b111100;
				8'b1000000: c <= 9'b101011000;
				8'b1110110: c <= 9'b100;
				8'b100101: c <= 9'b100000010;
				8'b101111: c <= 9'b11101100;
				8'b100110: c <= 9'b110001100;
				8'b1100011: c <= 9'b100110011;
				8'b1001000: c <= 9'b100101110;
				8'b111000: c <= 9'b10110100;
				8'b110001: c <= 9'b101010111;
				8'b1010111: c <= 9'b101010010;
				8'b1001110: c <= 9'b10000101;
				8'b1101010: c <= 9'b111010111;
				8'b1001001: c <= 9'b100010001;
				8'b1100000: c <= 9'b1111011;
				8'b110111: c <= 9'b100110111;
				8'b1011101: c <= 9'b111011111;
				8'b1011011: c <= 9'b110100101;
				8'b111001: c <= 9'b100011011;
				8'b1001010: c <= 9'b111000100;
				8'b110011: c <= 9'b110010111;
				8'b1101100: c <= 9'b11001100;
				8'b1110111: c <= 9'b101000010;
				8'b101011: c <= 9'b101111000;
				8'b1101011: c <= 9'b111001100;
				8'b111100: c <= 9'b110000000;
				8'b1000111: c <= 9'b10;
				8'b1011111: c <= 9'b11011001;
				8'b1110100: c <= 9'b1110111;
				8'b101101: c <= 9'b111000000;
				8'b1010011: c <= 9'b111011010;
				8'b1100001: c <= 9'b10110;
				8'b110101: c <= 9'b100111101;
				8'b1000100: c <= 9'b10001110;
				8'b1010001: c <= 9'b100001001;
				8'b1010100: c <= 9'b100100101;
				8'b1100110: c <= 9'b110110000;
				8'b101010: c <= 9'b111000111;
				8'b1011110: c <= 9'b101000001;
				8'b1100111: c <= 9'b10011;
				8'b1011010: c <= 9'b1111111;
				8'b1000010: c <= 9'b101101110;
				8'b111101: c <= 9'b110010001;
				8'b110000: c <= 9'b101000011;
				8'b111110: c <= 9'b100010011;
				8'b1100010: c <= 9'b101010111;
				8'b1110000: c <= 9'b11110011;
				8'b1101001: c <= 9'b1101010;
				8'b1110011: c <= 9'b111100011;
				8'b1001100: c <= 9'b111001101;
				8'b100001: c <= 9'b100011011;
				8'b1000110: c <= 9'b100110011;
				8'b1110010: c <= 9'b101100000;
				8'b1010000: c <= 9'b1101000;
				8'b1111010: c <= 9'b11001100;
				8'b1010101: c <= 9'b1111101;
				8'b111011: c <= 9'b111010001;
				8'b1001101: c <= 9'b101010000;
				8'b111111: c <= 9'b11001000;
				8'b1101110: c <= 9'b11000000;
				8'b1111011: c <= 9'b101010110;
				8'b1001011: c <= 9'b100110110;
				8'b1101111: c <= 9'b110101001;
				8'b1101000: c <= 9'b101000001;
				8'b101100: c <= 9'b100010;
				8'b100100: c <= 9'b1010101;
				8'b1111000: c <= 9'b100000000;
				8'b1000101: c <= 9'b101100000;
				8'b1011001: c <= 9'b100100011;
				8'b110100: c <= 9'b100000101;
				8'b1111001: c <= 9'b110101;
				8'b1110001: c <= 9'b111101101;
				8'b1001111: c <= 9'b111;
				8'b1100101: c <= 9'b111010010;
				8'b1111110: c <= 9'b110110010;
				8'b1111100: c <= 9'b1010000;
				8'b1010110: c <= 9'b111111;
				8'b110010: c <= 9'b101110011;
				8'b1101101: c <= 9'b11011001;
				8'b100011: c <= 9'b110001011;
				8'b1110101: c <= 9'b110111110;
				8'b1111101: c <= 9'b100000011;
				8'b101001: c <= 9'b100101001;
				8'b1010010: c <= 9'b101101001;
				8'b1011000: c <= 9'b100101110;
				8'b101110: c <= 9'b110110011;
				8'b1000001: c <= 9'b10111010;
				default: c <= 9'b0;
			endcase
			9'b111100 : case(di)
				8'b1000011: c <= 9'b1111000;
				8'b101000: c <= 9'b10000101;
				8'b111010: c <= 9'b100000110;
				8'b110110: c <= 9'b1001111;
				8'b1100100: c <= 9'b111101010;
				8'b1000000: c <= 9'b111100001;
				8'b1110110: c <= 9'b101010100;
				8'b100101: c <= 9'b1111001;
				8'b101111: c <= 9'b1000000;
				8'b100110: c <= 9'b110001101;
				8'b1100011: c <= 9'b1100000;
				8'b1001000: c <= 9'b101101001;
				8'b111000: c <= 9'b11001111;
				8'b110001: c <= 9'b111010000;
				8'b1010111: c <= 9'b100101010;
				8'b1001110: c <= 9'b11000100;
				8'b1101010: c <= 9'b10101101;
				8'b1001001: c <= 9'b110101011;
				8'b1100000: c <= 9'b101001010;
				8'b110111: c <= 9'b111101111;
				8'b1011101: c <= 9'b10111101;
				8'b1011011: c <= 9'b11111001;
				8'b111001: c <= 9'b100101000;
				8'b1001010: c <= 9'b110111001;
				8'b110011: c <= 9'b11101011;
				8'b1101100: c <= 9'b101;
				8'b1110111: c <= 9'b1001000;
				8'b101011: c <= 9'b1001100;
				8'b1101011: c <= 9'b11100111;
				8'b111100: c <= 9'b111101;
				8'b1000111: c <= 9'b10011100;
				8'b1011111: c <= 9'b100110111;
				8'b1110100: c <= 9'b111001101;
				8'b101101: c <= 9'b11100001;
				8'b1010011: c <= 9'b110001011;
				8'b1100001: c <= 9'b100111;
				8'b110101: c <= 9'b111100111;
				8'b1000100: c <= 9'b101101111;
				8'b1010001: c <= 9'b101000101;
				8'b1010100: c <= 9'b101111001;
				8'b1100110: c <= 9'b111101;
				8'b101010: c <= 9'b100000110;
				8'b1011110: c <= 9'b101011110;
				8'b1100111: c <= 9'b10111101;
				8'b1011010: c <= 9'b11011;
				8'b1000010: c <= 9'b11010101;
				8'b111101: c <= 9'b100111100;
				8'b110000: c <= 9'b11101000;
				8'b111110: c <= 9'b110001010;
				8'b1100010: c <= 9'b110101100;
				8'b1110000: c <= 9'b10000001;
				8'b1101001: c <= 9'b1100000;
				8'b1110011: c <= 9'b110000001;
				8'b1001100: c <= 9'b111111110;
				8'b100001: c <= 9'b1010010;
				8'b1000110: c <= 9'b11110101;
				8'b1110010: c <= 9'b10011001;
				8'b1010000: c <= 9'b11110010;
				8'b1111010: c <= 9'b101011101;
				8'b1010101: c <= 9'b101010110;
				8'b111011: c <= 9'b11110000;
				8'b1001101: c <= 9'b111010010;
				8'b111111: c <= 9'b110011111;
				8'b1101110: c <= 9'b101101011;
				8'b1111011: c <= 9'b11000011;
				8'b1001011: c <= 9'b100000010;
				8'b1101111: c <= 9'b10110010;
				8'b1101000: c <= 9'b111111011;
				8'b101100: c <= 9'b100010110;
				8'b100100: c <= 9'b110110;
				8'b1111000: c <= 9'b110111100;
				8'b1000101: c <= 9'b1001110;
				8'b1011001: c <= 9'b1110100;
				8'b110100: c <= 9'b110001010;
				8'b1111001: c <= 9'b110101110;
				8'b1110001: c <= 9'b1010111;
				8'b1001111: c <= 9'b111100001;
				8'b1100101: c <= 9'b101010001;
				8'b1111110: c <= 9'b111001;
				8'b1111100: c <= 9'b11111;
				8'b1010110: c <= 9'b110110;
				8'b110010: c <= 9'b10011100;
				8'b1101101: c <= 9'b100101101;
				8'b100011: c <= 9'b1011;
				8'b1110101: c <= 9'b101101110;
				8'b1111101: c <= 9'b100011000;
				8'b101001: c <= 9'b11011100;
				8'b1010010: c <= 9'b110000101;
				8'b1011000: c <= 9'b11101001;
				8'b101110: c <= 9'b110001101;
				8'b1000001: c <= 9'b11011001;
				default: c <= 9'b0;
			endcase
			9'b1010101 : case(di)
				8'b1000011: c <= 9'b110100001;
				8'b101000: c <= 9'b111101001;
				8'b111010: c <= 9'b11001101;
				8'b110110: c <= 9'b11101101;
				8'b1100100: c <= 9'b111111;
				8'b1000000: c <= 9'b111010010;
				8'b1110110: c <= 9'b101100101;
				8'b100101: c <= 9'b1011010;
				8'b101111: c <= 9'b110100000;
				8'b100110: c <= 9'b110011101;
				8'b1100011: c <= 9'b111010;
				8'b1001000: c <= 9'b10111011;
				8'b111000: c <= 9'b1100001;
				8'b110001: c <= 9'b101100100;
				8'b1010111: c <= 9'b10111011;
				8'b1001110: c <= 9'b101010101;
				8'b1101010: c <= 9'b1110010;
				8'b1001001: c <= 9'b1011110;
				8'b1100000: c <= 9'b110100000;
				8'b110111: c <= 9'b11111100;
				8'b1011101: c <= 9'b111101111;
				8'b1011011: c <= 9'b110110101;
				8'b111001: c <= 9'b10100000;
				8'b1001010: c <= 9'b11000100;
				8'b110011: c <= 9'b111001101;
				8'b1101100: c <= 9'b11111;
				8'b1110111: c <= 9'b10100010;
				8'b101011: c <= 9'b101000101;
				8'b1101011: c <= 9'b111000110;
				8'b111100: c <= 9'b101011001;
				8'b1000111: c <= 9'b101111000;
				8'b1011111: c <= 9'b100100000;
				8'b1110100: c <= 9'b101001;
				8'b101101: c <= 9'b110001010;
				8'b1010011: c <= 9'b100101010;
				8'b1100001: c <= 9'b11011101;
				8'b110101: c <= 9'b100100001;
				8'b1000100: c <= 9'b101010100;
				8'b1010001: c <= 9'b10010000;
				8'b1010100: c <= 9'b11110011;
				8'b1100110: c <= 9'b101010110;
				8'b101010: c <= 9'b11011001;
				8'b1011110: c <= 9'b11010111;
				8'b1100111: c <= 9'b1111;
				8'b1011010: c <= 9'b101000111;
				8'b1000010: c <= 9'b10110;
				8'b111101: c <= 9'b10001000;
				8'b110000: c <= 9'b111000011;
				8'b111110: c <= 9'b10110101;
				8'b1100010: c <= 9'b1011100;
				8'b1110000: c <= 9'b101011011;
				8'b1101001: c <= 9'b100001100;
				8'b1110011: c <= 9'b1010011;
				8'b1001100: c <= 9'b111;
				8'b100001: c <= 9'b100000001;
				8'b1000110: c <= 9'b101000100;
				8'b1110010: c <= 9'b111001;
				8'b1010000: c <= 9'b110111001;
				8'b1111010: c <= 9'b111000100;
				8'b1010101: c <= 9'b10010001;
				8'b111011: c <= 9'b111001010;
				8'b1001101: c <= 9'b110100010;
				8'b111111: c <= 9'b100111110;
				8'b1101110: c <= 9'b111111;
				8'b1111011: c <= 9'b10011111;
				8'b1001011: c <= 9'b10010111;
				8'b1101111: c <= 9'b10001000;
				8'b1101000: c <= 9'b1110100;
				8'b101100: c <= 9'b11111010;
				8'b100100: c <= 9'b100100;
				8'b1111000: c <= 9'b110001101;
				8'b1000101: c <= 9'b10001111;
				8'b1011001: c <= 9'b101010100;
				8'b110100: c <= 9'b100001110;
				8'b1111001: c <= 9'b100110110;
				8'b1110001: c <= 9'b11111000;
				8'b1001111: c <= 9'b1100111;
				8'b1100101: c <= 9'b110010110;
				8'b1111110: c <= 9'b110000101;
				8'b1111100: c <= 9'b11011000;
				8'b1010110: c <= 9'b10011;
				8'b110010: c <= 9'b1010001;
				8'b1101101: c <= 9'b10001100;
				8'b100011: c <= 9'b11011011;
				8'b1110101: c <= 9'b1111110;
				8'b1111101: c <= 9'b111000101;
				8'b101001: c <= 9'b101101000;
				8'b1010010: c <= 9'b111010111;
				8'b1011000: c <= 9'b10000;
				8'b101110: c <= 9'b110101;
				8'b1000001: c <= 9'b10110100;
				default: c <= 9'b0;
			endcase
			9'b11101111 : case(di)
				8'b1000011: c <= 9'b1110010;
				8'b101000: c <= 9'b10111110;
				8'b111010: c <= 9'b10100100;
				8'b110110: c <= 9'b100110010;
				8'b1100100: c <= 9'b10000111;
				8'b1000000: c <= 9'b111001101;
				8'b1110110: c <= 9'b10101101;
				8'b100101: c <= 9'b111101101;
				8'b101111: c <= 9'b111100010;
				8'b100110: c <= 9'b111000101;
				8'b1100011: c <= 9'b101110001;
				8'b1001000: c <= 9'b1111101;
				8'b111000: c <= 9'b10011011;
				8'b110001: c <= 9'b11100;
				8'b1010111: c <= 9'b100100101;
				8'b1001110: c <= 9'b110100100;
				8'b1101010: c <= 9'b100101011;
				8'b1001001: c <= 9'b101011101;
				8'b1100000: c <= 9'b111100000;
				8'b110111: c <= 9'b10100011;
				8'b1011101: c <= 9'b110011111;
				8'b1011011: c <= 9'b101011;
				8'b111001: c <= 9'b111110011;
				8'b1001010: c <= 9'b10100100;
				8'b110011: c <= 9'b11100010;
				8'b1101100: c <= 9'b110111111;
				8'b1110111: c <= 9'b11010010;
				8'b101011: c <= 9'b100011000;
				8'b1101011: c <= 9'b110010001;
				8'b111100: c <= 9'b1001111;
				8'b1000111: c <= 9'b1010110;
				8'b1011111: c <= 9'b101110110;
				8'b1110100: c <= 9'b1001111;
				8'b101101: c <= 9'b10101101;
				8'b1010011: c <= 9'b10111111;
				8'b1100001: c <= 9'b111011110;
				8'b110101: c <= 9'b100100001;
				8'b1000100: c <= 9'b101101110;
				8'b1010001: c <= 9'b100001111;
				8'b1010100: c <= 9'b111100100;
				8'b1100110: c <= 9'b100000011;
				8'b101010: c <= 9'b101101000;
				8'b1011110: c <= 9'b1001111;
				8'b1100111: c <= 9'b1000010;
				8'b1011010: c <= 9'b1101;
				8'b1000010: c <= 9'b11001111;
				8'b111101: c <= 9'b1111;
				8'b110000: c <= 9'b101001000;
				8'b111110: c <= 9'b10000110;
				8'b1100010: c <= 9'b100111011;
				8'b1110000: c <= 9'b110011010;
				8'b1101001: c <= 9'b1101101;
				8'b1110011: c <= 9'b1100001;
				8'b1001100: c <= 9'b1001;
				8'b100001: c <= 9'b111011011;
				8'b1000110: c <= 9'b100011;
				8'b1110010: c <= 9'b10101110;
				8'b1010000: c <= 9'b1101010;
				8'b1111010: c <= 9'b11010100;
				8'b1010101: c <= 9'b101110111;
				8'b111011: c <= 9'b1111011;
				8'b1001101: c <= 9'b10100111;
				8'b111111: c <= 9'b100010000;
				8'b1101110: c <= 9'b101110101;
				8'b1111011: c <= 9'b110100101;
				8'b1001011: c <= 9'b11000001;
				8'b1101111: c <= 9'b111101;
				8'b1101000: c <= 9'b111110110;
				8'b101100: c <= 9'b100001111;
				8'b100100: c <= 9'b110000001;
				8'b1111000: c <= 9'b111111110;
				8'b1000101: c <= 9'b101001011;
				8'b1011001: c <= 9'b1101010;
				8'b110100: c <= 9'b100000110;
				8'b1111001: c <= 9'b11110111;
				8'b1110001: c <= 9'b1001111;
				8'b1001111: c <= 9'b101100110;
				8'b1100101: c <= 9'b100000100;
				8'b1111110: c <= 9'b1101101;
				8'b1111100: c <= 9'b11111010;
				8'b1010110: c <= 9'b10001010;
				8'b110010: c <= 9'b111111011;
				8'b1101101: c <= 9'b10101101;
				8'b100011: c <= 9'b100011111;
				8'b1110101: c <= 9'b1111011;
				8'b1111101: c <= 9'b111101110;
				8'b101001: c <= 9'b11010001;
				8'b1010010: c <= 9'b110011;
				8'b1011000: c <= 9'b11111001;
				8'b101110: c <= 9'b110001110;
				8'b1000001: c <= 9'b10000111;
				default: c <= 9'b0;
			endcase
			9'b1011001 : case(di)
				8'b1000011: c <= 9'b110010111;
				8'b101000: c <= 9'b11101111;
				8'b111010: c <= 9'b1111011;
				8'b110110: c <= 9'b10100011;
				8'b1100100: c <= 9'b110100001;
				8'b1000000: c <= 9'b1011000;
				8'b1110110: c <= 9'b1000101;
				8'b100101: c <= 9'b110101111;
				8'b101111: c <= 9'b110001000;
				8'b100110: c <= 9'b111111001;
				8'b1100011: c <= 9'b100110111;
				8'b1001000: c <= 9'b101001110;
				8'b111000: c <= 9'b1111110;
				8'b110001: c <= 9'b101101101;
				8'b1010111: c <= 9'b111101;
				8'b1001110: c <= 9'b111101001;
				8'b1101010: c <= 9'b11010000;
				8'b1001001: c <= 9'b100100011;
				8'b1100000: c <= 9'b1111001;
				8'b110111: c <= 9'b101010101;
				8'b1011101: c <= 9'b101001100;
				8'b1011011: c <= 9'b11101101;
				8'b111001: c <= 9'b101000;
				8'b1001010: c <= 9'b101101001;
				8'b110011: c <= 9'b111101100;
				8'b1101100: c <= 9'b1110101;
				8'b1110111: c <= 9'b111011010;
				8'b101011: c <= 9'b11;
				8'b1101011: c <= 9'b10000101;
				8'b111100: c <= 9'b100110100;
				8'b1000111: c <= 9'b101000100;
				8'b1011111: c <= 9'b101011011;
				8'b1110100: c <= 9'b110101010;
				8'b101101: c <= 9'b1101111;
				8'b1010011: c <= 9'b11111110;
				8'b1100001: c <= 9'b10101101;
				8'b110101: c <= 9'b100001001;
				8'b1000100: c <= 9'b101111010;
				8'b1010001: c <= 9'b111100100;
				8'b1010100: c <= 9'b10000101;
				8'b1100110: c <= 9'b100110111;
				8'b101010: c <= 9'b110101111;
				8'b1011110: c <= 9'b100101100;
				8'b1100111: c <= 9'b10000010;
				8'b1011010: c <= 9'b111100001;
				8'b1000010: c <= 9'b11100100;
				8'b111101: c <= 9'b111101001;
				8'b110000: c <= 9'b110010100;
				8'b111110: c <= 9'b11110010;
				8'b1100010: c <= 9'b110100110;
				8'b1110000: c <= 9'b11001100;
				8'b1101001: c <= 9'b11100100;
				8'b1110011: c <= 9'b101110100;
				8'b1001100: c <= 9'b10001111;
				8'b100001: c <= 9'b100010011;
				8'b1000110: c <= 9'b11011010;
				8'b1110010: c <= 9'b1100;
				8'b1010000: c <= 9'b111101000;
				8'b1111010: c <= 9'b1101001;
				8'b1010101: c <= 9'b101110100;
				8'b111011: c <= 9'b101011000;
				8'b1001101: c <= 9'b110000011;
				8'b111111: c <= 9'b110011111;
				8'b1101110: c <= 9'b110011101;
				8'b1111011: c <= 9'b100111111;
				8'b1001011: c <= 9'b111010110;
				8'b1101111: c <= 9'b10111110;
				8'b1101000: c <= 9'b101100100;
				8'b101100: c <= 9'b11000111;
				8'b100100: c <= 9'b101100111;
				8'b1111000: c <= 9'b1101101;
				8'b1000101: c <= 9'b111101101;
				8'b1011001: c <= 9'b110111000;
				8'b110100: c <= 9'b111001101;
				8'b1111001: c <= 9'b111001010;
				8'b1110001: c <= 9'b10011101;
				8'b1001111: c <= 9'b110000101;
				8'b1100101: c <= 9'b1010000;
				8'b1111110: c <= 9'b100000011;
				8'b1111100: c <= 9'b110000;
				8'b1010110: c <= 9'b101101110;
				8'b110010: c <= 9'b1111000;
				8'b1101101: c <= 9'b111111110;
				8'b100011: c <= 9'b111111010;
				8'b1110101: c <= 9'b10010000;
				8'b1111101: c <= 9'b100101110;
				8'b101001: c <= 9'b10010111;
				8'b1010010: c <= 9'b100101001;
				8'b1011000: c <= 9'b101100101;
				8'b101110: c <= 9'b100001110;
				8'b1000001: c <= 9'b10000110;
				default: c <= 9'b0;
			endcase
			9'b11011011 : case(di)
				8'b1000011: c <= 9'b111111110;
				8'b101000: c <= 9'b11110000;
				8'b111010: c <= 9'b11110000;
				8'b110110: c <= 9'b10000111;
				8'b1100100: c <= 9'b101100;
				8'b1000000: c <= 9'b1110010;
				8'b1110110: c <= 9'b1111;
				8'b100101: c <= 9'b1110111;
				8'b101111: c <= 9'b10110100;
				8'b100110: c <= 9'b1000001;
				8'b1100011: c <= 9'b1001111;
				8'b1001000: c <= 9'b10010101;
				8'b111000: c <= 9'b11;
				8'b110001: c <= 9'b101100010;
				8'b1010111: c <= 9'b100000100;
				8'b1001110: c <= 9'b101110000;
				8'b1101010: c <= 9'b10010100;
				8'b1001001: c <= 9'b110101111;
				8'b1100000: c <= 9'b11100101;
				8'b110111: c <= 9'b100110110;
				8'b1011101: c <= 9'b110110110;
				8'b1011011: c <= 9'b110010101;
				8'b111001: c <= 9'b101010010;
				8'b1001010: c <= 9'b110001101;
				8'b110011: c <= 9'b110111010;
				8'b1101100: c <= 9'b101001100;
				8'b1110111: c <= 9'b11001110;
				8'b101011: c <= 9'b100010001;
				8'b1101011: c <= 9'b11001011;
				8'b111100: c <= 9'b100000000;
				8'b1000111: c <= 9'b10111110;
				8'b1011111: c <= 9'b11000110;
				8'b1110100: c <= 9'b1110;
				8'b101101: c <= 9'b101101011;
				8'b1010011: c <= 9'b100100101;
				8'b1100001: c <= 9'b11110110;
				8'b110101: c <= 9'b11001000;
				8'b1000100: c <= 9'b11100111;
				8'b1010001: c <= 9'b110000010;
				8'b1010100: c <= 9'b110111;
				8'b1100110: c <= 9'b10001001;
				8'b101010: c <= 9'b10011011;
				8'b1011110: c <= 9'b10001100;
				8'b1100111: c <= 9'b101010110;
				8'b1011010: c <= 9'b101010011;
				8'b1000010: c <= 9'b10111111;
				8'b111101: c <= 9'b110101110;
				8'b110000: c <= 9'b110101110;
				8'b111110: c <= 9'b1110010;
				8'b1100010: c <= 9'b1000000;
				8'b1110000: c <= 9'b11101;
				8'b1101001: c <= 9'b10010110;
				8'b1110011: c <= 9'b11111;
				8'b1001100: c <= 9'b10110011;
				8'b100001: c <= 9'b11010000;
				8'b1000110: c <= 9'b101001010;
				8'b1110010: c <= 9'b100110100;
				8'b1010000: c <= 9'b111010111;
				8'b1111010: c <= 9'b101101011;
				8'b1010101: c <= 9'b111101010;
				8'b111011: c <= 9'b11000111;
				8'b1001101: c <= 9'b1110010;
				8'b111111: c <= 9'b110110100;
				8'b1101110: c <= 9'b101001110;
				8'b1111011: c <= 9'b11010101;
				8'b1001011: c <= 9'b10110;
				8'b1101111: c <= 9'b111;
				8'b1101000: c <= 9'b11111010;
				8'b101100: c <= 9'b111100011;
				8'b100100: c <= 9'b10111000;
				8'b1111000: c <= 9'b11010111;
				8'b1000101: c <= 9'b101111111;
				8'b1011001: c <= 9'b1011011;
				8'b110100: c <= 9'b101000101;
				8'b1111001: c <= 9'b110011101;
				8'b1110001: c <= 9'b100100001;
				8'b1001111: c <= 9'b1101;
				8'b1100101: c <= 9'b110010001;
				8'b1111110: c <= 9'b1100100;
				8'b1111100: c <= 9'b1111101;
				8'b1010110: c <= 9'b101100100;
				8'b110010: c <= 9'b1011010;
				8'b1101101: c <= 9'b100111111;
				8'b100011: c <= 9'b1011100;
				8'b1110101: c <= 9'b111111110;
				8'b1111101: c <= 9'b110100;
				8'b101001: c <= 9'b1111111;
				8'b1010010: c <= 9'b10110;
				8'b1011000: c <= 9'b100011100;
				8'b101110: c <= 9'b110010101;
				8'b1000001: c <= 9'b110011011;
				default: c <= 9'b0;
			endcase
			9'b110001101 : case(di)
				8'b1000011: c <= 9'b10010101;
				8'b101000: c <= 9'b100011100;
				8'b111010: c <= 9'b100000111;
				8'b110110: c <= 9'b100000000;
				8'b1100100: c <= 9'b100001010;
				8'b1000000: c <= 9'b10111;
				8'b1110110: c <= 9'b101100011;
				8'b100101: c <= 9'b11010;
				8'b101111: c <= 9'b100000110;
				8'b100110: c <= 9'b110101101;
				8'b1100011: c <= 9'b10001001;
				8'b1001000: c <= 9'b101110101;
				8'b111000: c <= 9'b11001100;
				8'b110001: c <= 9'b111111;
				8'b1010111: c <= 9'b100100001;
				8'b1001110: c <= 9'b10111001;
				8'b1101010: c <= 9'b10000001;
				8'b1001001: c <= 9'b101001010;
				8'b1100000: c <= 9'b100100011;
				8'b110111: c <= 9'b111011011;
				8'b1011101: c <= 9'b1001001;
				8'b1011011: c <= 9'b10010001;
				8'b111001: c <= 9'b10010111;
				8'b1001010: c <= 9'b11001001;
				8'b110011: c <= 9'b10000011;
				8'b1101100: c <= 9'b11000010;
				8'b1110111: c <= 9'b111111;
				8'b101011: c <= 9'b100010111;
				8'b1101011: c <= 9'b1100100;
				8'b111100: c <= 9'b110111010;
				8'b1000111: c <= 9'b100001111;
				8'b1011111: c <= 9'b100000010;
				8'b1110100: c <= 9'b10101001;
				8'b101101: c <= 9'b101000110;
				8'b1010011: c <= 9'b111000100;
				8'b1100001: c <= 9'b111101010;
				8'b110101: c <= 9'b101010100;
				8'b1000100: c <= 9'b11001100;
				8'b1010001: c <= 9'b11110011;
				8'b1010100: c <= 9'b10000111;
				8'b1100110: c <= 9'b110000001;
				8'b101010: c <= 9'b100001011;
				8'b1011110: c <= 9'b110100100;
				8'b1100111: c <= 9'b111010;
				8'b1011010: c <= 9'b111101101;
				8'b1000010: c <= 9'b10110001;
				8'b111101: c <= 9'b111011;
				8'b110000: c <= 9'b11010000;
				8'b111110: c <= 9'b11111110;
				8'b1100010: c <= 9'b111101110;
				8'b1110000: c <= 9'b11000;
				8'b1101001: c <= 9'b11110100;
				8'b1110011: c <= 9'b111100010;
				8'b1001100: c <= 9'b11100110;
				8'b100001: c <= 9'b110000010;
				8'b1000110: c <= 9'b111100011;
				8'b1110010: c <= 9'b110000;
				8'b1010000: c <= 9'b111011100;
				8'b1111010: c <= 9'b100011001;
				8'b1010101: c <= 9'b1111010;
				8'b111011: c <= 9'b101011000;
				8'b1001101: c <= 9'b100111000;
				8'b111111: c <= 9'b100110000;
				8'b1101110: c <= 9'b11000011;
				8'b1111011: c <= 9'b111111010;
				8'b1001011: c <= 9'b110111000;
				8'b1101111: c <= 9'b101010000;
				8'b1101000: c <= 9'b1100100;
				8'b101100: c <= 9'b100011100;
				8'b100100: c <= 9'b111100000;
				8'b1111000: c <= 9'b101100010;
				8'b1000101: c <= 9'b11001111;
				8'b1011001: c <= 9'b11010;
				8'b110100: c <= 9'b101001011;
				8'b1111001: c <= 9'b100010101;
				8'b1110001: c <= 9'b100010010;
				8'b1001111: c <= 9'b10011011;
				8'b1100101: c <= 9'b10000010;
				8'b1111110: c <= 9'b10100;
				8'b1111100: c <= 9'b11101101;
				8'b1010110: c <= 9'b10111010;
				8'b110010: c <= 9'b111011111;
				8'b1101101: c <= 9'b10110110;
				8'b100011: c <= 9'b110100000;
				8'b1110101: c <= 9'b111100;
				8'b1111101: c <= 9'b1011001;
				8'b101001: c <= 9'b1101110;
				8'b1010010: c <= 9'b110111100;
				8'b1011000: c <= 9'b110100011;
				8'b101110: c <= 9'b101100110;
				8'b1000001: c <= 9'b110110;
				default: c <= 9'b0;
			endcase
			9'b11010011 : case(di)
				8'b1000011: c <= 9'b10010111;
				8'b101000: c <= 9'b101100101;
				8'b111010: c <= 9'b11001001;
				8'b110110: c <= 9'b10000010;
				8'b1100100: c <= 9'b11111011;
				8'b1000000: c <= 9'b11110011;
				8'b1110110: c <= 9'b101011011;
				8'b100101: c <= 9'b1010101;
				8'b101111: c <= 9'b100010;
				8'b100110: c <= 9'b110001001;
				8'b1100011: c <= 9'b1000;
				8'b1001000: c <= 9'b1010111;
				8'b111000: c <= 9'b100011111;
				8'b110001: c <= 9'b11011110;
				8'b1010111: c <= 9'b110110111;
				8'b1001110: c <= 9'b101101111;
				8'b1101010: c <= 9'b110010011;
				8'b1001001: c <= 9'b100001;
				8'b1100000: c <= 9'b101111000;
				8'b110111: c <= 9'b11111100;
				8'b1011101: c <= 9'b10000011;
				8'b1011011: c <= 9'b101011010;
				8'b111001: c <= 9'b1110000;
				8'b1001010: c <= 9'b101111001;
				8'b110011: c <= 9'b110010001;
				8'b1101100: c <= 9'b11001100;
				8'b1110111: c <= 9'b110101;
				8'b101011: c <= 9'b100101011;
				8'b1101011: c <= 9'b111011;
				8'b111100: c <= 9'b11001110;
				8'b1000111: c <= 9'b101000;
				8'b1011111: c <= 9'b111010000;
				8'b1110100: c <= 9'b11111000;
				8'b101101: c <= 9'b10011011;
				8'b1010011: c <= 9'b111101001;
				8'b1100001: c <= 9'b101100100;
				8'b110101: c <= 9'b101110010;
				8'b1000100: c <= 9'b110011110;
				8'b1010001: c <= 9'b11100100;
				8'b1010100: c <= 9'b110100111;
				8'b1100110: c <= 9'b110110100;
				8'b101010: c <= 9'b10011;
				8'b1011110: c <= 9'b1101;
				8'b1100111: c <= 9'b110101001;
				8'b1011010: c <= 9'b101101110;
				8'b1000010: c <= 9'b10100110;
				8'b111101: c <= 9'b111011;
				8'b110000: c <= 9'b111100010;
				8'b111110: c <= 9'b10011000;
				8'b1100010: c <= 9'b101011011;
				8'b1110000: c <= 9'b11010011;
				8'b1101001: c <= 9'b11110;
				8'b1110011: c <= 9'b101110110;
				8'b1001100: c <= 9'b100101;
				8'b100001: c <= 9'b110011110;
				8'b1000110: c <= 9'b10011;
				8'b1110010: c <= 9'b11101100;
				8'b1010000: c <= 9'b100111010;
				8'b1111010: c <= 9'b110010111;
				8'b1010101: c <= 9'b11111100;
				8'b111011: c <= 9'b111101010;
				8'b1001101: c <= 9'b100101;
				8'b111111: c <= 9'b10011101;
				8'b1101110: c <= 9'b111011010;
				8'b1111011: c <= 9'b110011111;
				8'b1001011: c <= 9'b100101000;
				8'b1101111: c <= 9'b111111;
				8'b1101000: c <= 9'b10111100;
				8'b101100: c <= 9'b1011100;
				8'b100100: c <= 9'b1110000;
				8'b1111000: c <= 9'b110010111;
				8'b1000101: c <= 9'b101110;
				8'b1011001: c <= 9'b111011101;
				8'b110100: c <= 9'b110011000;
				8'b1111001: c <= 9'b110001100;
				8'b1110001: c <= 9'b10000010;
				8'b1001111: c <= 9'b111111111;
				8'b1100101: c <= 9'b110000000;
				8'b1111110: c <= 9'b10001011;
				8'b1111100: c <= 9'b100000111;
				8'b1010110: c <= 9'b111001011;
				8'b110010: c <= 9'b11100000;
				8'b1101101: c <= 9'b110001100;
				8'b100011: c <= 9'b10000111;
				8'b1110101: c <= 9'b101101001;
				8'b1111101: c <= 9'b111010100;
				8'b101001: c <= 9'b101100110;
				8'b1010010: c <= 9'b10111;
				8'b1011000: c <= 9'b100000111;
				8'b101110: c <= 9'b11001011;
				8'b1000001: c <= 9'b1010111;
				default: c <= 9'b0;
			endcase
			9'b100010100 : case(di)
				8'b1000011: c <= 9'b10001100;
				8'b101000: c <= 9'b110111;
				8'b111010: c <= 9'b11000100;
				8'b110110: c <= 9'b101100000;
				8'b1100100: c <= 9'b10111110;
				8'b1000000: c <= 9'b10000110;
				8'b1110110: c <= 9'b1001000;
				8'b100101: c <= 9'b10010111;
				8'b101111: c <= 9'b101010111;
				8'b100110: c <= 9'b110001001;
				8'b1100011: c <= 9'b100101101;
				8'b1001000: c <= 9'b111101100;
				8'b111000: c <= 9'b111110110;
				8'b110001: c <= 9'b10010110;
				8'b1010111: c <= 9'b101000001;
				8'b1001110: c <= 9'b10110011;
				8'b1101010: c <= 9'b1001100;
				8'b1001001: c <= 9'b101101;
				8'b1100000: c <= 9'b110;
				8'b110111: c <= 9'b101011101;
				8'b1011101: c <= 9'b11010111;
				8'b1011011: c <= 9'b1001101;
				8'b111001: c <= 9'b100111111;
				8'b1001010: c <= 9'b111101001;
				8'b110011: c <= 9'b100111111;
				8'b1101100: c <= 9'b111101010;
				8'b1110111: c <= 9'b100010011;
				8'b101011: c <= 9'b100100000;
				8'b1101011: c <= 9'b1100100;
				8'b111100: c <= 9'b10011111;
				8'b1000111: c <= 9'b10111;
				8'b1011111: c <= 9'b1110001;
				8'b1110100: c <= 9'b1100010;
				8'b101101: c <= 9'b11010000;
				8'b1010011: c <= 9'b11010010;
				8'b1100001: c <= 9'b11111011;
				8'b110101: c <= 9'b100101110;
				8'b1000100: c <= 9'b10100010;
				8'b1010001: c <= 9'b101011101;
				8'b1010100: c <= 9'b100101001;
				8'b1100110: c <= 9'b10111001;
				8'b101010: c <= 9'b100110011;
				8'b1011110: c <= 9'b1101101;
				8'b1100111: c <= 9'b100111001;
				8'b1011010: c <= 9'b11111100;
				8'b1000010: c <= 9'b100011010;
				8'b111101: c <= 9'b110100011;
				8'b110000: c <= 9'b10010101;
				8'b111110: c <= 9'b1110101;
				8'b1100010: c <= 9'b1101000;
				8'b1110000: c <= 9'b101011000;
				8'b1101001: c <= 9'b111101000;
				8'b1110011: c <= 9'b110100000;
				8'b1001100: c <= 9'b10010111;
				8'b100001: c <= 9'b111011110;
				8'b1000110: c <= 9'b111100110;
				8'b1110010: c <= 9'b10111001;
				8'b1010000: c <= 9'b111111110;
				8'b1111010: c <= 9'b1101101;
				8'b1010101: c <= 9'b100100001;
				8'b111011: c <= 9'b101010;
				8'b1001101: c <= 9'b10100;
				8'b111111: c <= 9'b10110101;
				8'b1101110: c <= 9'b100000110;
				8'b1111011: c <= 9'b100101010;
				8'b1001011: c <= 9'b100011100;
				8'b1101111: c <= 9'b111001011;
				8'b1101000: c <= 9'b1101010;
				8'b101100: c <= 9'b11101001;
				8'b100100: c <= 9'b100001;
				8'b1111000: c <= 9'b111000110;
				8'b1000101: c <= 9'b11000011;
				8'b1011001: c <= 9'b11100100;
				8'b110100: c <= 9'b100100101;
				8'b1111001: c <= 9'b1100001;
				8'b1110001: c <= 9'b1001101;
				8'b1001111: c <= 9'b110000;
				8'b1100101: c <= 9'b111110000;
				8'b1111110: c <= 9'b10000110;
				8'b1111100: c <= 9'b111011101;
				8'b1010110: c <= 9'b11110000;
				8'b110010: c <= 9'b100001;
				8'b1101101: c <= 9'b110101011;
				8'b100011: c <= 9'b100011010;
				8'b1110101: c <= 9'b100111001;
				8'b1111101: c <= 9'b110001100;
				8'b101001: c <= 9'b1101010;
				8'b1010010: c <= 9'b1110;
				8'b1011000: c <= 9'b111010100;
				8'b101110: c <= 9'b1000000;
				8'b1000001: c <= 9'b110011110;
				default: c <= 9'b0;
			endcase
			9'b101101 : case(di)
				8'b1000011: c <= 9'b111010110;
				8'b101000: c <= 9'b110100101;
				8'b111010: c <= 9'b111000110;
				8'b110110: c <= 9'b110010010;
				8'b1100100: c <= 9'b110000111;
				8'b1000000: c <= 9'b110110101;
				8'b1110110: c <= 9'b111000111;
				8'b100101: c <= 9'b11;
				8'b101111: c <= 9'b101101110;
				8'b100110: c <= 9'b110110100;
				8'b1100011: c <= 9'b10011100;
				8'b1001000: c <= 9'b1101101;
				8'b111000: c <= 9'b10111010;
				8'b110001: c <= 9'b11010101;
				8'b1010111: c <= 9'b11111010;
				8'b1001110: c <= 9'b101011110;
				8'b1101010: c <= 9'b11110;
				8'b1001001: c <= 9'b1101101;
				8'b1100000: c <= 9'b100010111;
				8'b110111: c <= 9'b101101011;
				8'b1011101: c <= 9'b111100101;
				8'b1011011: c <= 9'b10101011;
				8'b111001: c <= 9'b10001100;
				8'b1001010: c <= 9'b110111010;
				8'b110011: c <= 9'b1110;
				8'b1101100: c <= 9'b100110100;
				8'b1110111: c <= 9'b1;
				8'b101011: c <= 9'b1010111;
				8'b1101011: c <= 9'b101110010;
				8'b111100: c <= 9'b111111011;
				8'b1000111: c <= 9'b110100101;
				8'b1011111: c <= 9'b11101100;
				8'b1110100: c <= 9'b11110110;
				8'b101101: c <= 9'b1001100;
				8'b1010011: c <= 9'b111111010;
				8'b1100001: c <= 9'b111101001;
				8'b110101: c <= 9'b10101011;
				8'b1000100: c <= 9'b10111100;
				8'b1010001: c <= 9'b100101001;
				8'b1010100: c <= 9'b101100100;
				8'b1100110: c <= 9'b10001001;
				8'b101010: c <= 9'b11110011;
				8'b1011110: c <= 9'b101000001;
				8'b1100111: c <= 9'b1011100;
				8'b1011010: c <= 9'b100010100;
				8'b1000010: c <= 9'b1000010;
				8'b111101: c <= 9'b10101010;
				8'b110000: c <= 9'b110101111;
				8'b111110: c <= 9'b1011011;
				8'b1100010: c <= 9'b111100011;
				8'b1110000: c <= 9'b11100001;
				8'b1101001: c <= 9'b111010;
				8'b1110011: c <= 9'b10101010;
				8'b1001100: c <= 9'b1111010;
				8'b100001: c <= 9'b110100000;
				8'b1000110: c <= 9'b10110001;
				8'b1110010: c <= 9'b11010100;
				8'b1010000: c <= 9'b10101100;
				8'b1111010: c <= 9'b1111000;
				8'b1010101: c <= 9'b11110101;
				8'b111011: c <= 9'b101101101;
				8'b1001101: c <= 9'b1011100;
				8'b111111: c <= 9'b100000000;
				8'b1101110: c <= 9'b100010010;
				8'b1111011: c <= 9'b100001111;
				8'b1001011: c <= 9'b1110000;
				8'b1101111: c <= 9'b11010000;
				8'b1101000: c <= 9'b111010111;
				8'b101100: c <= 9'b101110011;
				8'b100100: c <= 9'b11001010;
				8'b1111000: c <= 9'b10010001;
				8'b1000101: c <= 9'b11100;
				8'b1011001: c <= 9'b1111001;
				8'b110100: c <= 9'b1100010;
				8'b1111001: c <= 9'b100000110;
				8'b1110001: c <= 9'b100011;
				8'b1001111: c <= 9'b111010100;
				8'b1100101: c <= 9'b111100001;
				8'b1111110: c <= 9'b100001;
				8'b1111100: c <= 9'b1111110;
				8'b1010110: c <= 9'b110100001;
				8'b110010: c <= 9'b100001001;
				8'b1101101: c <= 9'b11010101;
				8'b100011: c <= 9'b100011101;
				8'b1110101: c <= 9'b100010100;
				8'b1111101: c <= 9'b11010100;
				8'b101001: c <= 9'b10001010;
				8'b1010010: c <= 9'b11010100;
				8'b1011000: c <= 9'b11100;
				8'b101110: c <= 9'b10011011;
				8'b1000001: c <= 9'b10110001;
				default: c <= 9'b0;
			endcase
			9'b10101010 : case(di)
				8'b1000011: c <= 9'b11111001;
				8'b101000: c <= 9'b11001100;
				8'b111010: c <= 9'b110101011;
				8'b110110: c <= 9'b101110001;
				8'b1100100: c <= 9'b110110011;
				8'b1000000: c <= 9'b10101101;
				8'b1110110: c <= 9'b111011101;
				8'b100101: c <= 9'b110000001;
				8'b101111: c <= 9'b1001100;
				8'b100110: c <= 9'b101011010;
				8'b1100011: c <= 9'b111100011;
				8'b1001000: c <= 9'b111100001;
				8'b111000: c <= 9'b101101;
				8'b110001: c <= 9'b101110110;
				8'b1010111: c <= 9'b100101010;
				8'b1001110: c <= 9'b111011010;
				8'b1101010: c <= 9'b110010011;
				8'b1001001: c <= 9'b1111;
				8'b1100000: c <= 9'b1101100;
				8'b110111: c <= 9'b100101100;
				8'b1011101: c <= 9'b101;
				8'b1011011: c <= 9'b101001110;
				8'b111001: c <= 9'b1000000;
				8'b1001010: c <= 9'b111111101;
				8'b110011: c <= 9'b110100111;
				8'b1101100: c <= 9'b100101001;
				8'b1110111: c <= 9'b11110111;
				8'b101011: c <= 9'b111011100;
				8'b1101011: c <= 9'b101100100;
				8'b111100: c <= 9'b10000010;
				8'b1000111: c <= 9'b100000010;
				8'b1011111: c <= 9'b101100;
				8'b1110100: c <= 9'b111010100;
				8'b101101: c <= 9'b100101110;
				8'b1010011: c <= 9'b111100100;
				8'b1100001: c <= 9'b111101000;
				8'b110101: c <= 9'b10011000;
				8'b1000100: c <= 9'b10010001;
				8'b1010001: c <= 9'b11111000;
				8'b1010100: c <= 9'b1011000;
				8'b1100110: c <= 9'b10010000;
				8'b101010: c <= 9'b10010110;
				8'b1011110: c <= 9'b10001010;
				8'b1100111: c <= 9'b101001011;
				8'b1011010: c <= 9'b110111;
				8'b1000010: c <= 9'b100011101;
				8'b111101: c <= 9'b11001100;
				8'b110000: c <= 9'b101010000;
				8'b111110: c <= 9'b11011;
				8'b1100010: c <= 9'b100000100;
				8'b1110000: c <= 9'b101100101;
				8'b1101001: c <= 9'b101110010;
				8'b1110011: c <= 9'b110111000;
				8'b1001100: c <= 9'b101;
				8'b100001: c <= 9'b110011;
				8'b1000110: c <= 9'b11110101;
				8'b1110010: c <= 9'b110100111;
				8'b1010000: c <= 9'b10101111;
				8'b1111010: c <= 9'b10101111;
				8'b1010101: c <= 9'b111011110;
				8'b111011: c <= 9'b100000100;
				8'b1001101: c <= 9'b111110110;
				8'b111111: c <= 9'b110111010;
				8'b1101110: c <= 9'b110001;
				8'b1111011: c <= 9'b100001010;
				8'b1001011: c <= 9'b101011111;
				8'b1101111: c <= 9'b1010110;
				8'b1101000: c <= 9'b10010100;
				8'b101100: c <= 9'b10111;
				8'b100100: c <= 9'b111101;
				8'b1111000: c <= 9'b111100111;
				8'b1000101: c <= 9'b11001011;
				8'b1011001: c <= 9'b101110001;
				8'b110100: c <= 9'b111101010;
				8'b1111001: c <= 9'b1000111;
				8'b1110001: c <= 9'b101000001;
				8'b1001111: c <= 9'b11110;
				8'b1100101: c <= 9'b110100100;
				8'b1111110: c <= 9'b11111010;
				8'b1111100: c <= 9'b10110100;
				8'b1010110: c <= 9'b111101010;
				8'b110010: c <= 9'b1000111;
				8'b1101101: c <= 9'b100111111;
				8'b100011: c <= 9'b101100111;
				8'b1110101: c <= 9'b101101;
				8'b1111101: c <= 9'b111111010;
				8'b101001: c <= 9'b100100110;
				8'b1010010: c <= 9'b1100001;
				8'b1011000: c <= 9'b100101;
				8'b101110: c <= 9'b111010;
				8'b1000001: c <= 9'b100011010;
				default: c <= 9'b0;
			endcase
			9'b11111 : case(di)
				8'b1000011: c <= 9'b1010011;
				8'b101000: c <= 9'b111111000;
				8'b111010: c <= 9'b1101101;
				8'b110110: c <= 9'b111001;
				8'b1100100: c <= 9'b10001010;
				8'b1000000: c <= 9'b11011000;
				8'b1110110: c <= 9'b111110000;
				8'b100101: c <= 9'b1100011;
				8'b101111: c <= 9'b111101;
				8'b100110: c <= 9'b111001001;
				8'b1100011: c <= 9'b111011100;
				8'b1001000: c <= 9'b10001010;
				8'b111000: c <= 9'b100010110;
				8'b110001: c <= 9'b100100010;
				8'b1010111: c <= 9'b11100;
				8'b1001110: c <= 9'b100101100;
				8'b1101010: c <= 9'b10;
				8'b1001001: c <= 9'b10111110;
				8'b1100000: c <= 9'b100101001;
				8'b110111: c <= 9'b1000110;
				8'b1011101: c <= 9'b111101101;
				8'b1011011: c <= 9'b101100010;
				8'b111001: c <= 9'b101010;
				8'b1001010: c <= 9'b1101001;
				8'b110011: c <= 9'b10001110;
				8'b1101100: c <= 9'b100101000;
				8'b1110111: c <= 9'b110110111;
				8'b101011: c <= 9'b100000111;
				8'b1101011: c <= 9'b101110010;
				8'b111100: c <= 9'b10110101;
				8'b1000111: c <= 9'b110001100;
				8'b1011111: c <= 9'b10111011;
				8'b1110100: c <= 9'b11000000;
				8'b101101: c <= 9'b101101000;
				8'b1010011: c <= 9'b100111110;
				8'b1100001: c <= 9'b110100;
				8'b110101: c <= 9'b110101011;
				8'b1000100: c <= 9'b110100010;
				8'b1010001: c <= 9'b110011001;
				8'b1010100: c <= 9'b111001010;
				8'b1100110: c <= 9'b1011011;
				8'b101010: c <= 9'b1000;
				8'b1011110: c <= 9'b11000111;
				8'b1100111: c <= 9'b101011001;
				8'b1011010: c <= 9'b1110;
				8'b1000010: c <= 9'b100100010;
				8'b111101: c <= 9'b1100;
				8'b110000: c <= 9'b111101101;
				8'b111110: c <= 9'b11110010;
				8'b1100010: c <= 9'b111101101;
				8'b1110000: c <= 9'b100011010;
				8'b1101001: c <= 9'b10110011;
				8'b1110011: c <= 9'b101110100;
				8'b1001100: c <= 9'b100111111;
				8'b100001: c <= 9'b1101001;
				8'b1000110: c <= 9'b110011;
				8'b1110010: c <= 9'b10111111;
				8'b1010000: c <= 9'b110100000;
				8'b1111010: c <= 9'b100011000;
				8'b1010101: c <= 9'b110111010;
				8'b111011: c <= 9'b1111011;
				8'b1001101: c <= 9'b110010010;
				8'b111111: c <= 9'b110011;
				8'b1101110: c <= 9'b111111010;
				8'b1111011: c <= 9'b101101011;
				8'b1001011: c <= 9'b111001111;
				8'b1101111: c <= 9'b1001011;
				8'b1101000: c <= 9'b1010010;
				8'b101100: c <= 9'b100000000;
				8'b100100: c <= 9'b11101011;
				8'b1111000: c <= 9'b10111011;
				8'b1000101: c <= 9'b110011001;
				8'b1011001: c <= 9'b1000101;
				8'b110100: c <= 9'b101110010;
				8'b1111001: c <= 9'b1010011;
				8'b1110001: c <= 9'b111101101;
				8'b1001111: c <= 9'b111000;
				8'b1100101: c <= 9'b110101110;
				8'b1111110: c <= 9'b11011011;
				8'b1111100: c <= 9'b101101110;
				8'b1010110: c <= 9'b110000011;
				8'b110010: c <= 9'b11010011;
				8'b1101101: c <= 9'b1110001;
				8'b100011: c <= 9'b110000001;
				8'b1110101: c <= 9'b101000111;
				8'b1111101: c <= 9'b100000101;
				8'b101001: c <= 9'b110101110;
				8'b1010010: c <= 9'b101000001;
				8'b1011000: c <= 9'b110110011;
				8'b101110: c <= 9'b11010011;
				8'b1000001: c <= 9'b1101101;
				default: c <= 9'b0;
			endcase
			9'b100001001 : case(di)
				8'b1000011: c <= 9'b11100000;
				8'b101000: c <= 9'b101101111;
				8'b111010: c <= 9'b1001100;
				8'b110110: c <= 9'b101011111;
				8'b1100100: c <= 9'b11100001;
				8'b1000000: c <= 9'b100100111;
				8'b1110110: c <= 9'b101011010;
				8'b100101: c <= 9'b101010;
				8'b101111: c <= 9'b11100;
				8'b100110: c <= 9'b110010111;
				8'b1100011: c <= 9'b1001;
				8'b1001000: c <= 9'b1001100;
				8'b111000: c <= 9'b1011011;
				8'b110001: c <= 9'b100011000;
				8'b1010111: c <= 9'b110101010;
				8'b1001110: c <= 9'b111001;
				8'b1101010: c <= 9'b100001010;
				8'b1001001: c <= 9'b111001110;
				8'b1100000: c <= 9'b101011000;
				8'b110111: c <= 9'b10;
				8'b1011101: c <= 9'b110001101;
				8'b1011011: c <= 9'b101100001;
				8'b111001: c <= 9'b100100001;
				8'b1001010: c <= 9'b101100011;
				8'b110011: c <= 9'b10001010;
				8'b1101100: c <= 9'b100100111;
				8'b1110111: c <= 9'b10011111;
				8'b101011: c <= 9'b11011;
				8'b1101011: c <= 9'b111000000;
				8'b111100: c <= 9'b100001011;
				8'b1000111: c <= 9'b101000100;
				8'b1011111: c <= 9'b111111110;
				8'b1110100: c <= 9'b11011000;
				8'b101101: c <= 9'b100110111;
				8'b1010011: c <= 9'b11111011;
				8'b1100001: c <= 9'b110001100;
				8'b110101: c <= 9'b111101100;
				8'b1000100: c <= 9'b111110001;
				8'b1010001: c <= 9'b100101101;
				8'b1010100: c <= 9'b101101100;
				8'b1100110: c <= 9'b100101011;
				8'b101010: c <= 9'b1001001;
				8'b1011110: c <= 9'b1110111;
				8'b1100111: c <= 9'b11111;
				8'b1011010: c <= 9'b110101;
				8'b1000010: c <= 9'b1100010;
				8'b111101: c <= 9'b1001000;
				8'b110000: c <= 9'b110011101;
				8'b111110: c <= 9'b11100000;
				8'b1100010: c <= 9'b111101001;
				8'b1110000: c <= 9'b100001010;
				8'b1101001: c <= 9'b110011100;
				8'b1110011: c <= 9'b11110100;
				8'b1001100: c <= 9'b101111001;
				8'b100001: c <= 9'b110001;
				8'b1000110: c <= 9'b101100;
				8'b1110010: c <= 9'b100010110;
				8'b1010000: c <= 9'b1011011;
				8'b1111010: c <= 9'b11000011;
				8'b1010101: c <= 9'b101011111;
				8'b111011: c <= 9'b100010011;
				8'b1001101: c <= 9'b10101110;
				8'b111111: c <= 9'b10001110;
				8'b1101110: c <= 9'b10001011;
				8'b1111011: c <= 9'b100000100;
				8'b1001011: c <= 9'b101110010;
				8'b1101111: c <= 9'b10110111;
				8'b1101000: c <= 9'b101101000;
				8'b101100: c <= 9'b110001101;
				8'b100100: c <= 9'b1110011;
				8'b1111000: c <= 9'b1110100;
				8'b1000101: c <= 9'b11000010;
				8'b1011001: c <= 9'b110;
				8'b110100: c <= 9'b100111;
				8'b1111001: c <= 9'b10101;
				8'b1110001: c <= 9'b1000001;
				8'b1001111: c <= 9'b100100011;
				8'b1100101: c <= 9'b1100010;
				8'b1111110: c <= 9'b1001100;
				8'b1111100: c <= 9'b101010000;
				8'b1010110: c <= 9'b111011110;
				8'b110010: c <= 9'b100110011;
				8'b1101101: c <= 9'b100010011;
				8'b100011: c <= 9'b1000110;
				8'b1110101: c <= 9'b1000;
				8'b1111101: c <= 9'b111110101;
				8'b101001: c <= 9'b111100100;
				8'b1010010: c <= 9'b11011100;
				8'b1011000: c <= 9'b1001101;
				8'b101110: c <= 9'b1100001;
				8'b1000001: c <= 9'b1100010;
				default: c <= 9'b0;
			endcase
			9'b101101000 : case(di)
				8'b1000011: c <= 9'b101001100;
				8'b101000: c <= 9'b10101001;
				8'b111010: c <= 9'b110010001;
				8'b110110: c <= 9'b111001100;
				8'b1100100: c <= 9'b111001101;
				8'b1000000: c <= 9'b110000010;
				8'b1110110: c <= 9'b101111010;
				8'b100101: c <= 9'b1100110;
				8'b101111: c <= 9'b1111000;
				8'b100110: c <= 9'b10110110;
				8'b1100011: c <= 9'b101101000;
				8'b1001000: c <= 9'b1000001;
				8'b111000: c <= 9'b100110010;
				8'b110001: c <= 9'b100101110;
				8'b1010111: c <= 9'b10011010;
				8'b1001110: c <= 9'b11101101;
				8'b1101010: c <= 9'b110100100;
				8'b1001001: c <= 9'b1000000;
				8'b1100000: c <= 9'b111011111;
				8'b110111: c <= 9'b1011011;
				8'b1011101: c <= 9'b11000111;
				8'b1011011: c <= 9'b1010110;
				8'b111001: c <= 9'b1001100;
				8'b1001010: c <= 9'b1101101;
				8'b110011: c <= 9'b10100100;
				8'b1101100: c <= 9'b10110100;
				8'b1110111: c <= 9'b110001011;
				8'b101011: c <= 9'b10010111;
				8'b1101011: c <= 9'b101101;
				8'b111100: c <= 9'b101100111;
				8'b1000111: c <= 9'b110100001;
				8'b1011111: c <= 9'b11101100;
				8'b1110100: c <= 9'b1110000;
				8'b101101: c <= 9'b10101001;
				8'b1010011: c <= 9'b100111;
				8'b1100001: c <= 9'b1001110;
				8'b110101: c <= 9'b101011000;
				8'b1000100: c <= 9'b11111011;
				8'b1010001: c <= 9'b1001000;
				8'b1010100: c <= 9'b111111;
				8'b1100110: c <= 9'b10000010;
				8'b101010: c <= 9'b110110011;
				8'b1011110: c <= 9'b11111110;
				8'b1100111: c <= 9'b111111000;
				8'b1011010: c <= 9'b100000001;
				8'b1000010: c <= 9'b10011;
				8'b111101: c <= 9'b111011111;
				8'b110000: c <= 9'b10101100;
				8'b111110: c <= 9'b110000;
				8'b1100010: c <= 9'b11000111;
				8'b1110000: c <= 9'b11010010;
				8'b1101001: c <= 9'b11011011;
				8'b1110011: c <= 9'b100100101;
				8'b1001100: c <= 9'b10000010;
				8'b100001: c <= 9'b1000;
				8'b1000110: c <= 9'b100110;
				8'b1110010: c <= 9'b110011101;
				8'b1010000: c <= 9'b101101;
				8'b1111010: c <= 9'b101111001;
				8'b1010101: c <= 9'b100010011;
				8'b111011: c <= 9'b100111110;
				8'b1001101: c <= 9'b1111010;
				8'b111111: c <= 9'b101011111;
				8'b1101110: c <= 9'b100111001;
				8'b1111011: c <= 9'b111010;
				8'b1001011: c <= 9'b110000110;
				8'b1101111: c <= 9'b1100100;
				8'b1101000: c <= 9'b1100010;
				8'b101100: c <= 9'b101111110;
				8'b100100: c <= 9'b1111;
				8'b1111000: c <= 9'b110001111;
				8'b1000101: c <= 9'b111110011;
				8'b1011001: c <= 9'b11100100;
				8'b110100: c <= 9'b101100001;
				8'b1111001: c <= 9'b110010010;
				8'b1110001: c <= 9'b100100110;
				8'b1001111: c <= 9'b11010100;
				8'b1100101: c <= 9'b10110110;
				8'b1111110: c <= 9'b101111000;
				8'b1111100: c <= 9'b111001000;
				8'b1010110: c <= 9'b100011111;
				8'b110010: c <= 9'b101001010;
				8'b1101101: c <= 9'b11111101;
				8'b100011: c <= 9'b100111;
				8'b1110101: c <= 9'b110100001;
				8'b1111101: c <= 9'b11110011;
				8'b101001: c <= 9'b10001001;
				8'b1010010: c <= 9'b110001100;
				8'b1011000: c <= 9'b1111000;
				8'b101110: c <= 9'b11000;
				8'b1000001: c <= 9'b11100111;
				default: c <= 9'b0;
			endcase
			9'b11111001 : case(di)
				8'b1000011: c <= 9'b1100001;
				8'b101000: c <= 9'b101110000;
				8'b111010: c <= 9'b101011110;
				8'b110110: c <= 9'b110001100;
				8'b1100100: c <= 9'b111010110;
				8'b1000000: c <= 9'b1110100;
				8'b1110110: c <= 9'b110011000;
				8'b100101: c <= 9'b1011111;
				8'b101111: c <= 9'b100010101;
				8'b100110: c <= 9'b10000101;
				8'b1100011: c <= 9'b111011001;
				8'b1001000: c <= 9'b11010111;
				8'b111000: c <= 9'b111100011;
				8'b110001: c <= 9'b110011010;
				8'b1010111: c <= 9'b100000110;
				8'b1001110: c <= 9'b110000101;
				8'b1101010: c <= 9'b1101010;
				8'b1001001: c <= 9'b10101101;
				8'b1100000: c <= 9'b100011111;
				8'b110111: c <= 9'b111111000;
				8'b1011101: c <= 9'b110001001;
				8'b1011011: c <= 9'b100111000;
				8'b111001: c <= 9'b111001001;
				8'b1001010: c <= 9'b11101000;
				8'b110011: c <= 9'b10010001;
				8'b1101100: c <= 9'b100001101;
				8'b1110111: c <= 9'b10101101;
				8'b101011: c <= 9'b101110100;
				8'b1101011: c <= 9'b100000101;
				8'b111100: c <= 9'b101010001;
				8'b1000111: c <= 9'b10101110;
				8'b1011111: c <= 9'b100100001;
				8'b1110100: c <= 9'b111000100;
				8'b101101: c <= 9'b11011010;
				8'b1010011: c <= 9'b11101;
				8'b1100001: c <= 9'b100001001;
				8'b110101: c <= 9'b111011010;
				8'b1000100: c <= 9'b1;
				8'b1010001: c <= 9'b101110000;
				8'b1010100: c <= 9'b100010;
				8'b1100110: c <= 9'b1001110;
				8'b101010: c <= 9'b1110001;
				8'b1011110: c <= 9'b100010110;
				8'b1100111: c <= 9'b111000110;
				8'b1011010: c <= 9'b101001111;
				8'b1000010: c <= 9'b101110010;
				8'b111101: c <= 9'b110001000;
				8'b110000: c <= 9'b100000110;
				8'b111110: c <= 9'b101010101;
				8'b1100010: c <= 9'b110101100;
				8'b1110000: c <= 9'b100110100;
				8'b1101001: c <= 9'b10101010;
				8'b1110011: c <= 9'b110111111;
				8'b1001100: c <= 9'b111111010;
				8'b100001: c <= 9'b101011111;
				8'b1000110: c <= 9'b11101101;
				8'b1110010: c <= 9'b100101101;
				8'b1010000: c <= 9'b10111010;
				8'b1111010: c <= 9'b110011010;
				8'b1010101: c <= 9'b10;
				8'b111011: c <= 9'b11110;
				8'b1001101: c <= 9'b11111000;
				8'b111111: c <= 9'b10000001;
				8'b1101110: c <= 9'b10011;
				8'b1111011: c <= 9'b11;
				8'b1001011: c <= 9'b10000001;
				8'b1101111: c <= 9'b110001101;
				8'b1101000: c <= 9'b100101000;
				8'b101100: c <= 9'b100010010;
				8'b100100: c <= 9'b11001011;
				8'b1111000: c <= 9'b110011010;
				8'b1000101: c <= 9'b10001110;
				8'b1011001: c <= 9'b1001111;
				8'b110100: c <= 9'b110000011;
				8'b1111001: c <= 9'b111001000;
				8'b1110001: c <= 9'b100111000;
				8'b1001111: c <= 9'b11010011;
				8'b1100101: c <= 9'b100101000;
				8'b1111110: c <= 9'b110000010;
				8'b1111100: c <= 9'b11100111;
				8'b1010110: c <= 9'b11111010;
				8'b110010: c <= 9'b110110000;
				8'b1101101: c <= 9'b10100101;
				8'b100011: c <= 9'b110010100;
				8'b1110101: c <= 9'b111000110;
				8'b1111101: c <= 9'b100100001;
				8'b101001: c <= 9'b101000111;
				8'b1010010: c <= 9'b111100100;
				8'b1011000: c <= 9'b100111111;
				8'b101110: c <= 9'b111101110;
				8'b1000001: c <= 9'b1011010;
				default: c <= 9'b0;
			endcase
			9'b11111110 : case(di)
				8'b1000011: c <= 9'b110011;
				8'b101000: c <= 9'b1001001;
				8'b111010: c <= 9'b1110;
				8'b110110: c <= 9'b10100011;
				8'b1100100: c <= 9'b111001001;
				8'b1000000: c <= 9'b111101110;
				8'b1110110: c <= 9'b1001001;
				8'b100101: c <= 9'b111101100;
				8'b101111: c <= 9'b1110101;
				8'b100110: c <= 9'b111001010;
				8'b1100011: c <= 9'b1000101;
				8'b1001000: c <= 9'b10001101;
				8'b111000: c <= 9'b1110001;
				8'b110001: c <= 9'b10111101;
				8'b1010111: c <= 9'b110111000;
				8'b1001110: c <= 9'b101100011;
				8'b1101010: c <= 9'b100110110;
				8'b1001001: c <= 9'b110000000;
				8'b1100000: c <= 9'b101011001;
				8'b110111: c <= 9'b1001010;
				8'b1011101: c <= 9'b111100011;
				8'b1011011: c <= 9'b110101;
				8'b111001: c <= 9'b110011000;
				8'b1001010: c <= 9'b101000100;
				8'b110011: c <= 9'b11100001;
				8'b1101100: c <= 9'b10010110;
				8'b1110111: c <= 9'b11001001;
				8'b101011: c <= 9'b100110010;
				8'b1101011: c <= 9'b101111010;
				8'b111100: c <= 9'b100101011;
				8'b1000111: c <= 9'b11001111;
				8'b1011111: c <= 9'b111101;
				8'b1110100: c <= 9'b1011110;
				8'b101101: c <= 9'b11010100;
				8'b1010011: c <= 9'b110011;
				8'b1100001: c <= 9'b11011101;
				8'b110101: c <= 9'b111111;
				8'b1000100: c <= 9'b110101010;
				8'b1010001: c <= 9'b101001000;
				8'b1010100: c <= 9'b100110101;
				8'b1100110: c <= 9'b111100010;
				8'b101010: c <= 9'b111010000;
				8'b1011110: c <= 9'b110101100;
				8'b1100111: c <= 9'b10001000;
				8'b1011010: c <= 9'b111;
				8'b1000010: c <= 9'b1010001;
				8'b111101: c <= 9'b100101000;
				8'b110000: c <= 9'b11001000;
				8'b111110: c <= 9'b11000100;
				8'b1100010: c <= 9'b100111000;
				8'b1110000: c <= 9'b11000110;
				8'b1101001: c <= 9'b110110000;
				8'b1110011: c <= 9'b11001101;
				8'b1001100: c <= 9'b100111100;
				8'b100001: c <= 9'b10111;
				8'b1000110: c <= 9'b111111000;
				8'b1110010: c <= 9'b100110010;
				8'b1010000: c <= 9'b100110010;
				8'b1111010: c <= 9'b10011001;
				8'b1010101: c <= 9'b100011;
				8'b111011: c <= 9'b10010101;
				8'b1001101: c <= 9'b100011;
				8'b111111: c <= 9'b101101101;
				8'b1101110: c <= 9'b1000101;
				8'b1111011: c <= 9'b110100011;
				8'b1001011: c <= 9'b110011000;
				8'b1101111: c <= 9'b110010110;
				8'b1101000: c <= 9'b100100001;
				8'b101100: c <= 9'b100;
				8'b100100: c <= 9'b1101110;
				8'b1111000: c <= 9'b11100011;
				8'b1000101: c <= 9'b1100111;
				8'b1011001: c <= 9'b110100101;
				8'b110100: c <= 9'b110111111;
				8'b1111001: c <= 9'b10001010;
				8'b1110001: c <= 9'b10100;
				8'b1001111: c <= 9'b100101110;
				8'b1100101: c <= 9'b11101;
				8'b1111110: c <= 9'b10010001;
				8'b1111100: c <= 9'b10011001;
				8'b1010110: c <= 9'b111010111;
				8'b110010: c <= 9'b111111101;
				8'b1101101: c <= 9'b101010111;
				8'b100011: c <= 9'b1100000;
				8'b1110101: c <= 9'b110011010;
				8'b1111101: c <= 9'b1000100;
				8'b101001: c <= 9'b110011001;
				8'b1010010: c <= 9'b100100001;
				8'b1011000: c <= 9'b11011;
				8'b101110: c <= 9'b111111011;
				8'b1000001: c <= 9'b101000011;
				default: c <= 9'b0;
			endcase
			9'b10110 : case(di)
				8'b1000011: c <= 9'b110101111;
				8'b101000: c <= 9'b1110011;
				8'b111010: c <= 9'b100000010;
				8'b110110: c <= 9'b10011;
				8'b1100100: c <= 9'b101010;
				8'b1000000: c <= 9'b1110001;
				8'b1110110: c <= 9'b111110001;
				8'b100101: c <= 9'b101101001;
				8'b101111: c <= 9'b111101001;
				8'b100110: c <= 9'b11000000;
				8'b1100011: c <= 9'b100110111;
				8'b1001000: c <= 9'b101101011;
				8'b111000: c <= 9'b101001010;
				8'b110001: c <= 9'b11101001;
				8'b1010111: c <= 9'b1011100;
				8'b1001110: c <= 9'b100101111;
				8'b1101010: c <= 9'b100111101;
				8'b1001001: c <= 9'b110110000;
				8'b1100000: c <= 9'b1110010;
				8'b110111: c <= 9'b101001100;
				8'b1011101: c <= 9'b101000111;
				8'b1011011: c <= 9'b111010111;
				8'b111001: c <= 9'b100010111;
				8'b1001010: c <= 9'b110010010;
				8'b110011: c <= 9'b110000010;
				8'b1101100: c <= 9'b111000;
				8'b1110111: c <= 9'b10101000;
				8'b101011: c <= 9'b110111111;
				8'b1101011: c <= 9'b111010000;
				8'b111100: c <= 9'b101101000;
				8'b1000111: c <= 9'b110011000;
				8'b1011111: c <= 9'b110001101;
				8'b1110100: c <= 9'b101110011;
				8'b101101: c <= 9'b100110;
				8'b1010011: c <= 9'b111011;
				8'b1100001: c <= 9'b101101001;
				8'b110101: c <= 9'b111100001;
				8'b1000100: c <= 9'b10110010;
				8'b1010001: c <= 9'b11011011;
				8'b1010100: c <= 9'b1111010;
				8'b1100110: c <= 9'b100100;
				8'b101010: c <= 9'b11100000;
				8'b1011110: c <= 9'b111111010;
				8'b1100111: c <= 9'b100001;
				8'b1011010: c <= 9'b10010;
				8'b1000010: c <= 9'b110000010;
				8'b111101: c <= 9'b111000000;
				8'b110000: c <= 9'b100101110;
				8'b111110: c <= 9'b11;
				8'b1100010: c <= 9'b100000100;
				8'b1110000: c <= 9'b11011000;
				8'b1101001: c <= 9'b1101101;
				8'b1110011: c <= 9'b111001;
				8'b1001100: c <= 9'b101110;
				8'b100001: c <= 9'b100001;
				8'b1000110: c <= 9'b1001110;
				8'b1110010: c <= 9'b110100111;
				8'b1010000: c <= 9'b110101010;
				8'b1111010: c <= 9'b111000111;
				8'b1010101: c <= 9'b10100111;
				8'b111011: c <= 9'b11010111;
				8'b1001101: c <= 9'b111110000;
				8'b111111: c <= 9'b10101100;
				8'b1101110: c <= 9'b100001010;
				8'b1111011: c <= 9'b111011011;
				8'b1001011: c <= 9'b100110;
				8'b1101111: c <= 9'b110000010;
				8'b1101000: c <= 9'b1111111;
				8'b101100: c <= 9'b11110001;
				8'b100100: c <= 9'b110001100;
				8'b1111000: c <= 9'b110100;
				8'b1000101: c <= 9'b10010111;
				8'b1011001: c <= 9'b11011000;
				8'b110100: c <= 9'b100101;
				8'b1111001: c <= 9'b1001100;
				8'b1110001: c <= 9'b1010001;
				8'b1001111: c <= 9'b11000111;
				8'b1100101: c <= 9'b1010101;
				8'b1111110: c <= 9'b100000111;
				8'b1111100: c <= 9'b1101001;
				8'b1010110: c <= 9'b11100101;
				8'b110010: c <= 9'b10011111;
				8'b1101101: c <= 9'b101110100;
				8'b100011: c <= 9'b111111;
				8'b1110101: c <= 9'b1110010;
				8'b1111101: c <= 9'b100111111;
				8'b101001: c <= 9'b10010000;
				8'b1010010: c <= 9'b10001011;
				8'b1011000: c <= 9'b1100111;
				8'b101110: c <= 9'b11111110;
				8'b1000001: c <= 9'b10010011;
				default: c <= 9'b0;
			endcase
			9'b101000111 : case(di)
				8'b1000011: c <= 9'b11111100;
				8'b101000: c <= 9'b111000111;
				8'b111010: c <= 9'b101111111;
				8'b110110: c <= 9'b110010100;
				8'b1100100: c <= 9'b100011101;
				8'b1000000: c <= 9'b11110001;
				8'b1110110: c <= 9'b100000101;
				8'b100101: c <= 9'b101010;
				8'b101111: c <= 9'b110101101;
				8'b100110: c <= 9'b11001101;
				8'b1100011: c <= 9'b110011001;
				8'b1001000: c <= 9'b100110100;
				8'b111000: c <= 9'b111000011;
				8'b110001: c <= 9'b11100000;
				8'b1010111: c <= 9'b1000001;
				8'b1001110: c <= 9'b100001111;
				8'b1101010: c <= 9'b100110111;
				8'b1001001: c <= 9'b1101;
				8'b1100000: c <= 9'b110011011;
				8'b110111: c <= 9'b10010;
				8'b1011101: c <= 9'b101000101;
				8'b1011011: c <= 9'b110100011;
				8'b111001: c <= 9'b101001100;
				8'b1001010: c <= 9'b100011011;
				8'b110011: c <= 9'b10100010;
				8'b1101100: c <= 9'b1101110;
				8'b1110111: c <= 9'b101001000;
				8'b101011: c <= 9'b10001000;
				8'b1101011: c <= 9'b10011001;
				8'b111100: c <= 9'b100100011;
				8'b1000111: c <= 9'b1;
				8'b1011111: c <= 9'b101110000;
				8'b1110100: c <= 9'b100111;
				8'b101101: c <= 9'b10000111;
				8'b1010011: c <= 9'b11;
				8'b1100001: c <= 9'b101000101;
				8'b110101: c <= 9'b10110110;
				8'b1000100: c <= 9'b110110;
				8'b1010001: c <= 9'b10001010;
				8'b1010100: c <= 9'b10011101;
				8'b1100110: c <= 9'b111001101;
				8'b101010: c <= 9'b111111001;
				8'b1011110: c <= 9'b101100000;
				8'b1100111: c <= 9'b1001011;
				8'b1011010: c <= 9'b101100011;
				8'b1000010: c <= 9'b101;
				8'b111101: c <= 9'b10011011;
				8'b110000: c <= 9'b11000110;
				8'b111110: c <= 9'b11010001;
				8'b1100010: c <= 9'b111100100;
				8'b1110000: c <= 9'b10110111;
				8'b1101001: c <= 9'b100101011;
				8'b1110011: c <= 9'b110100001;
				8'b1001100: c <= 9'b11010001;
				8'b100001: c <= 9'b110000001;
				8'b1000110: c <= 9'b10110010;
				8'b1110010: c <= 9'b10011011;
				8'b1010000: c <= 9'b10010101;
				8'b1111010: c <= 9'b101011000;
				8'b1010101: c <= 9'b11011010;
				8'b111011: c <= 9'b11000111;
				8'b1001101: c <= 9'b1000000;
				8'b111111: c <= 9'b10100;
				8'b1101110: c <= 9'b1001110;
				8'b1111011: c <= 9'b100100;
				8'b1001011: c <= 9'b101000001;
				8'b1101111: c <= 9'b11100110;
				8'b1101000: c <= 9'b10011;
				8'b101100: c <= 9'b101101111;
				8'b100100: c <= 9'b100111000;
				8'b1111000: c <= 9'b100101010;
				8'b1000101: c <= 9'b101011111;
				8'b1011001: c <= 9'b110001;
				8'b110100: c <= 9'b10000001;
				8'b1111001: c <= 9'b100010011;
				8'b1110001: c <= 9'b111110011;
				8'b1001111: c <= 9'b100101011;
				8'b1100101: c <= 9'b11101001;
				8'b1111110: c <= 9'b101101110;
				8'b1111100: c <= 9'b11110000;
				8'b1010110: c <= 9'b110001111;
				8'b110010: c <= 9'b101110;
				8'b1101101: c <= 9'b111011;
				8'b100011: c <= 9'b11110111;
				8'b1110101: c <= 9'b10100000;
				8'b1111101: c <= 9'b100111101;
				8'b101001: c <= 9'b111101101;
				8'b1010010: c <= 9'b1011100;
				8'b1011000: c <= 9'b110110;
				8'b101110: c <= 9'b110010001;
				8'b1000001: c <= 9'b111101001;
				default: c <= 9'b0;
			endcase
			9'b110100110 : case(di)
				8'b1000011: c <= 9'b100011100;
				8'b101000: c <= 9'b10000101;
				8'b111010: c <= 9'b11010001;
				8'b110110: c <= 9'b100111010;
				8'b1100100: c <= 9'b1110;
				8'b1000000: c <= 9'b1100010;
				8'b1110110: c <= 9'b110101111;
				8'b100101: c <= 9'b100100110;
				8'b101111: c <= 9'b111100110;
				8'b100110: c <= 9'b101000110;
				8'b1100011: c <= 9'b101001011;
				8'b1001000: c <= 9'b11110111;
				8'b111000: c <= 9'b101110100;
				8'b110001: c <= 9'b110100111;
				8'b1010111: c <= 9'b101010;
				8'b1001110: c <= 9'b1101100;
				8'b1101010: c <= 9'b100011000;
				8'b1001001: c <= 9'b10010110;
				8'b1100000: c <= 9'b1001111;
				8'b110111: c <= 9'b111010010;
				8'b1011101: c <= 9'b111001110;
				8'b1011011: c <= 9'b11000010;
				8'b111001: c <= 9'b11001111;
				8'b1001010: c <= 9'b101001;
				8'b110011: c <= 9'b100101;
				8'b1101100: c <= 9'b100100011;
				8'b1110111: c <= 9'b101101010;
				8'b101011: c <= 9'b1110111;
				8'b1101011: c <= 9'b101110;
				8'b111100: c <= 9'b110000110;
				8'b1000111: c <= 9'b100101011;
				8'b1011111: c <= 9'b10100111;
				8'b1110100: c <= 9'b100;
				8'b101101: c <= 9'b101101011;
				8'b1010011: c <= 9'b101111000;
				8'b1100001: c <= 9'b100111110;
				8'b110101: c <= 9'b111101000;
				8'b1000100: c <= 9'b1101000;
				8'b1010001: c <= 9'b100010;
				8'b1010100: c <= 9'b1011001;
				8'b1100110: c <= 9'b101001010;
				8'b101010: c <= 9'b1010110;
				8'b1011110: c <= 9'b10010;
				8'b1100111: c <= 9'b111101;
				8'b1011010: c <= 9'b11110000;
				8'b1000010: c <= 9'b100010011;
				8'b111101: c <= 9'b10101111;
				8'b110000: c <= 9'b110101110;
				8'b111110: c <= 9'b10100100;
				8'b1100010: c <= 9'b110110110;
				8'b1110000: c <= 9'b1101000;
				8'b1101001: c <= 9'b11011100;
				8'b1110011: c <= 9'b1100110;
				8'b1001100: c <= 9'b11110001;
				8'b100001: c <= 9'b1010010;
				8'b1000110: c <= 9'b111101;
				8'b1110010: c <= 9'b110010;
				8'b1010000: c <= 9'b1001111;
				8'b1111010: c <= 9'b100110011;
				8'b1010101: c <= 9'b11011110;
				8'b111011: c <= 9'b111010010;
				8'b1001101: c <= 9'b10010101;
				8'b111111: c <= 9'b11100111;
				8'b1101110: c <= 9'b1011000;
				8'b1111011: c <= 9'b11000111;
				8'b1001011: c <= 9'b100110000;
				8'b1101111: c <= 9'b10011100;
				8'b1101000: c <= 9'b10011001;
				8'b101100: c <= 9'b10101100;
				8'b100100: c <= 9'b100101101;
				8'b1111000: c <= 9'b100010100;
				8'b1000101: c <= 9'b11011011;
				8'b1011001: c <= 9'b101000110;
				8'b110100: c <= 9'b100011001;
				8'b1111001: c <= 9'b11100001;
				8'b1110001: c <= 9'b100000111;
				8'b1001111: c <= 9'b11011011;
				8'b1100101: c <= 9'b11011001;
				8'b1111110: c <= 9'b110001001;
				8'b1111100: c <= 9'b100100001;
				8'b1010110: c <= 9'b101101001;
				8'b110010: c <= 9'b100011001;
				8'b1101101: c <= 9'b1100000;
				8'b100011: c <= 9'b1000010;
				8'b1110101: c <= 9'b10110101;
				8'b1111101: c <= 9'b11001011;
				8'b101001: c <= 9'b101010010;
				8'b1010010: c <= 9'b101100010;
				8'b1011000: c <= 9'b110111010;
				8'b101110: c <= 9'b11011110;
				8'b1000001: c <= 9'b1101110;
				default: c <= 9'b0;
			endcase
			9'b111001101 : case(di)
				8'b1000011: c <= 9'b10010110;
				8'b101000: c <= 9'b101001011;
				8'b111010: c <= 9'b110010001;
				8'b110110: c <= 9'b100001111;
				8'b1100100: c <= 9'b111001110;
				8'b1000000: c <= 9'b1100101;
				8'b1110110: c <= 9'b11100001;
				8'b100101: c <= 9'b10100110;
				8'b101111: c <= 9'b110001101;
				8'b100110: c <= 9'b111001111;
				8'b1100011: c <= 9'b10101101;
				8'b1001000: c <= 9'b100100110;
				8'b111000: c <= 9'b10011010;
				8'b110001: c <= 9'b110000111;
				8'b1010111: c <= 9'b10100100;
				8'b1001110: c <= 9'b1010010;
				8'b1101010: c <= 9'b1111001;
				8'b1001001: c <= 9'b111000011;
				8'b1100000: c <= 9'b10100;
				8'b110111: c <= 9'b11100010;
				8'b1011101: c <= 9'b111001111;
				8'b1011011: c <= 9'b100111111;
				8'b111001: c <= 9'b10100011;
				8'b1001010: c <= 9'b11111001;
				8'b110011: c <= 9'b100010110;
				8'b1101100: c <= 9'b11110100;
				8'b1110111: c <= 9'b100111101;
				8'b101011: c <= 9'b110110110;
				8'b1101011: c <= 9'b11000001;
				8'b111100: c <= 9'b10100000;
				8'b1000111: c <= 9'b111100100;
				8'b1011111: c <= 9'b10001100;
				8'b1110100: c <= 9'b11011100;
				8'b101101: c <= 9'b111011110;
				8'b1010011: c <= 9'b10001111;
				8'b1100001: c <= 9'b101001110;
				8'b110101: c <= 9'b100110100;
				8'b1000100: c <= 9'b11111010;
				8'b1010001: c <= 9'b11111000;
				8'b1010100: c <= 9'b111001100;
				8'b1100110: c <= 9'b110011101;
				8'b101010: c <= 9'b111100101;
				8'b1011110: c <= 9'b1100110;
				8'b1100111: c <= 9'b110011111;
				8'b1011010: c <= 9'b111101111;
				8'b1000010: c <= 9'b110001111;
				8'b111101: c <= 9'b1010101;
				8'b110000: c <= 9'b101010101;
				8'b111110: c <= 9'b110111;
				8'b1100010: c <= 9'b111001101;
				8'b1110000: c <= 9'b11101000;
				8'b1101001: c <= 9'b100100110;
				8'b1110011: c <= 9'b1011001;
				8'b1001100: c <= 9'b10100110;
				8'b100001: c <= 9'b110111110;
				8'b1000110: c <= 9'b101010111;
				8'b1110010: c <= 9'b1111;
				8'b1010000: c <= 9'b10110101;
				8'b1111010: c <= 9'b101101000;
				8'b1010101: c <= 9'b1001111;
				8'b111011: c <= 9'b11011011;
				8'b1001101: c <= 9'b11010111;
				8'b111111: c <= 9'b100010010;
				8'b1101110: c <= 9'b100000001;
				8'b1111011: c <= 9'b100101;
				8'b1001011: c <= 9'b1101110;
				8'b1101111: c <= 9'b10000;
				8'b1101000: c <= 9'b111001101;
				8'b101100: c <= 9'b111000111;
				8'b100100: c <= 9'b101011001;
				8'b1111000: c <= 9'b1000101;
				8'b1000101: c <= 9'b111000110;
				8'b1011001: c <= 9'b1010101;
				8'b110100: c <= 9'b111010100;
				8'b1111001: c <= 9'b101111110;
				8'b1110001: c <= 9'b1011011;
				8'b1001111: c <= 9'b100101101;
				8'b1100101: c <= 9'b110101101;
				8'b1111110: c <= 9'b10110110;
				8'b1111100: c <= 9'b100100110;
				8'b1010110: c <= 9'b101101111;
				8'b110010: c <= 9'b10010110;
				8'b1101101: c <= 9'b111101111;
				8'b100011: c <= 9'b111111101;
				8'b1110101: c <= 9'b10110011;
				8'b1111101: c <= 9'b1001100;
				8'b101001: c <= 9'b110000010;
				8'b1010010: c <= 9'b110101011;
				8'b1011000: c <= 9'b101010000;
				8'b101110: c <= 9'b10111100;
				8'b1000001: c <= 9'b1000;
				default: c <= 9'b0;
			endcase
			9'b111101 : case(di)
				8'b1000011: c <= 9'b11101000;
				8'b101000: c <= 9'b100111;
				8'b111010: c <= 9'b1000001;
				8'b110110: c <= 9'b110100100;
				8'b1100100: c <= 9'b100101;
				8'b1000000: c <= 9'b110100101;
				8'b1110110: c <= 9'b101101110;
				8'b100101: c <= 9'b10111110;
				8'b101111: c <= 9'b101000100;
				8'b100110: c <= 9'b111001101;
				8'b1100011: c <= 9'b110000111;
				8'b1001000: c <= 9'b1000110;
				8'b111000: c <= 9'b11111;
				8'b110001: c <= 9'b1111000;
				8'b1010111: c <= 9'b11;
				8'b1001110: c <= 9'b10100000;
				8'b1101010: c <= 9'b100100;
				8'b1001001: c <= 9'b111011010;
				8'b1100000: c <= 9'b111000100;
				8'b110111: c <= 9'b10101101;
				8'b1011101: c <= 9'b100011000;
				8'b1011011: c <= 9'b10101101;
				8'b111001: c <= 9'b111010000;
				8'b1001010: c <= 9'b110100;
				8'b110011: c <= 9'b10110001;
				8'b1101100: c <= 9'b11011101;
				8'b1110111: c <= 9'b110000011;
				8'b101011: c <= 9'b101010110;
				8'b1101011: c <= 9'b100001111;
				8'b111100: c <= 9'b1101001;
				8'b1000111: c <= 9'b10110011;
				8'b1011111: c <= 9'b111111101;
				8'b1110100: c <= 9'b110101010;
				8'b101101: c <= 9'b10110110;
				8'b1010011: c <= 9'b11110100;
				8'b1100001: c <= 9'b110101011;
				8'b110101: c <= 9'b10011;
				8'b1000100: c <= 9'b110101001;
				8'b1010001: c <= 9'b111001011;
				8'b1010100: c <= 9'b111110000;
				8'b1100110: c <= 9'b11100001;
				8'b101010: c <= 9'b1001100;
				8'b1011110: c <= 9'b11010000;
				8'b1100111: c <= 9'b100010010;
				8'b1011010: c <= 9'b1111011;
				8'b1000010: c <= 9'b11001;
				8'b111101: c <= 9'b100110;
				8'b110000: c <= 9'b10110111;
				8'b111110: c <= 9'b100011100;
				8'b1100010: c <= 9'b101100110;
				8'b1110000: c <= 9'b10000001;
				8'b1101001: c <= 9'b10110001;
				8'b1110011: c <= 9'b1110001;
				8'b1001100: c <= 9'b11011101;
				8'b100001: c <= 9'b11001010;
				8'b1000110: c <= 9'b100111010;
				8'b1110010: c <= 9'b10101;
				8'b1010000: c <= 9'b101010111;
				8'b1111010: c <= 9'b101010;
				8'b1010101: c <= 9'b11101001;
				8'b111011: c <= 9'b1001011;
				8'b1001101: c <= 9'b1001100;
				8'b111111: c <= 9'b10101010;
				8'b1101110: c <= 9'b100100001;
				8'b1111011: c <= 9'b110011001;
				8'b1001011: c <= 9'b10100110;
				8'b1101111: c <= 9'b11011110;
				8'b1101000: c <= 9'b101000011;
				8'b101100: c <= 9'b10000;
				8'b100100: c <= 9'b110101011;
				8'b1111000: c <= 9'b100101100;
				8'b1000101: c <= 9'b100011100;
				8'b1011001: c <= 9'b1;
				8'b110100: c <= 9'b10100101;
				8'b1111001: c <= 9'b11011110;
				8'b1110001: c <= 9'b110001000;
				8'b1001111: c <= 9'b100110000;
				8'b1100101: c <= 9'b1001011;
				8'b1111110: c <= 9'b10110110;
				8'b1111100: c <= 9'b11010010;
				8'b1010110: c <= 9'b10101011;
				8'b110010: c <= 9'b100110011;
				8'b1101101: c <= 9'b11110111;
				8'b100011: c <= 9'b10001110;
				8'b1110101: c <= 9'b101100000;
				8'b1111101: c <= 9'b10001000;
				8'b101001: c <= 9'b100000010;
				8'b1010010: c <= 9'b10101001;
				8'b1011000: c <= 9'b11111010;
				8'b101110: c <= 9'b111111010;
				8'b1000001: c <= 9'b101101011;
				default: c <= 9'b0;
			endcase
			9'b110000101 : case(di)
				8'b1000011: c <= 9'b101001000;
				8'b101000: c <= 9'b110000110;
				8'b111010: c <= 9'b10001110;
				8'b110110: c <= 9'b1100011;
				8'b1100100: c <= 9'b110000;
				8'b1000000: c <= 9'b11000001;
				8'b1110110: c <= 9'b101111000;
				8'b100101: c <= 9'b100001010;
				8'b101111: c <= 9'b100100001;
				8'b100110: c <= 9'b101001100;
				8'b1100011: c <= 9'b1111101;
				8'b1001000: c <= 9'b11010001;
				8'b111000: c <= 9'b100110;
				8'b110001: c <= 9'b101101111;
				8'b1010111: c <= 9'b10000001;
				8'b1001110: c <= 9'b11111101;
				8'b1101010: c <= 9'b10110001;
				8'b1001001: c <= 9'b110101001;
				8'b1100000: c <= 9'b100010001;
				8'b110111: c <= 9'b110011001;
				8'b1011101: c <= 9'b101000010;
				8'b1011011: c <= 9'b101111000;
				8'b111001: c <= 9'b110100011;
				8'b1001010: c <= 9'b11011;
				8'b110011: c <= 9'b10111011;
				8'b1101100: c <= 9'b1010000;
				8'b1110111: c <= 9'b111010001;
				8'b101011: c <= 9'b110000011;
				8'b1101011: c <= 9'b11001111;
				8'b111100: c <= 9'b10111111;
				8'b1000111: c <= 9'b111011010;
				8'b1011111: c <= 9'b10100010;
				8'b1110100: c <= 9'b101101010;
				8'b101101: c <= 9'b100010;
				8'b1010011: c <= 9'b11011011;
				8'b1100001: c <= 9'b100010011;
				8'b110101: c <= 9'b10100111;
				8'b1000100: c <= 9'b10000;
				8'b1010001: c <= 9'b10101110;
				8'b1010100: c <= 9'b1101;
				8'b1100110: c <= 9'b110000111;
				8'b101010: c <= 9'b11011110;
				8'b1011110: c <= 9'b1101101;
				8'b1100111: c <= 9'b111111110;
				8'b1011010: c <= 9'b1101101;
				8'b1000010: c <= 9'b111101111;
				8'b111101: c <= 9'b1110000;
				8'b110000: c <= 9'b10111011;
				8'b111110: c <= 9'b101100001;
				8'b1100010: c <= 9'b1111100;
				8'b1110000: c <= 9'b101101101;
				8'b1101001: c <= 9'b100111100;
				8'b1110011: c <= 9'b101001010;
				8'b1001100: c <= 9'b101000011;
				8'b100001: c <= 9'b11000001;
				8'b1000110: c <= 9'b101100101;
				8'b1110010: c <= 9'b10010000;
				8'b1010000: c <= 9'b100101100;
				8'b1111010: c <= 9'b11000110;
				8'b1010101: c <= 9'b100111;
				8'b111011: c <= 9'b11100;
				8'b1001101: c <= 9'b111100011;
				8'b111111: c <= 9'b1001011;
				8'b1101110: c <= 9'b111100000;
				8'b1111011: c <= 9'b10101010;
				8'b1001011: c <= 9'b111111;
				8'b1101111: c <= 9'b100010101;
				8'b1101000: c <= 9'b101100101;
				8'b101100: c <= 9'b100011111;
				8'b100100: c <= 9'b11101111;
				8'b1111000: c <= 9'b11110110;
				8'b1000101: c <= 9'b110010101;
				8'b1011001: c <= 9'b101011110;
				8'b110100: c <= 9'b110000;
				8'b1111001: c <= 9'b110010110;
				8'b1110001: c <= 9'b101101;
				8'b1001111: c <= 9'b111010000;
				8'b1100101: c <= 9'b100100010;
				8'b1111110: c <= 9'b11000110;
				8'b1111100: c <= 9'b1100111;
				8'b1010110: c <= 9'b101010100;
				8'b110010: c <= 9'b101110011;
				8'b1101101: c <= 9'b10010011;
				8'b100011: c <= 9'b11100010;
				8'b1110101: c <= 9'b111011;
				8'b1111101: c <= 9'b10000101;
				8'b101001: c <= 9'b111001110;
				8'b1010010: c <= 9'b110110;
				8'b1011000: c <= 9'b10100011;
				8'b101110: c <= 9'b10011101;
				8'b1000001: c <= 9'b110;
				default: c <= 9'b0;
			endcase
			9'b1110010 : case(di)
				8'b1000011: c <= 9'b11001110;
				8'b101000: c <= 9'b1111110;
				8'b111010: c <= 9'b111100111;
				8'b110110: c <= 9'b110010100;
				8'b1100100: c <= 9'b110001010;
				8'b1000000: c <= 9'b100111001;
				8'b1110110: c <= 9'b111101100;
				8'b100101: c <= 9'b110101111;
				8'b101111: c <= 9'b1111010;
				8'b100110: c <= 9'b110000010;
				8'b1100011: c <= 9'b101000100;
				8'b1001000: c <= 9'b110101101;
				8'b111000: c <= 9'b101101000;
				8'b110001: c <= 9'b100101011;
				8'b1010111: c <= 9'b111100000;
				8'b1001110: c <= 9'b100101100;
				8'b1101010: c <= 9'b11010100;
				8'b1001001: c <= 9'b11001;
				8'b1100000: c <= 9'b111111111;
				8'b110111: c <= 9'b110011;
				8'b1011101: c <= 9'b11001101;
				8'b1011011: c <= 9'b111001001;
				8'b111001: c <= 9'b110010111;
				8'b1001010: c <= 9'b10010111;
				8'b110011: c <= 9'b110001011;
				8'b1101100: c <= 9'b101001011;
				8'b1110111: c <= 9'b1101101;
				8'b101011: c <= 9'b110101111;
				8'b1101011: c <= 9'b10111101;
				8'b111100: c <= 9'b1000100;
				8'b1000111: c <= 9'b10111101;
				8'b1011111: c <= 9'b10110110;
				8'b1110100: c <= 9'b110000111;
				8'b101101: c <= 9'b10001010;
				8'b1010011: c <= 9'b100000011;
				8'b1100001: c <= 9'b11100111;
				8'b110101: c <= 9'b11111011;
				8'b1000100: c <= 9'b1000011;
				8'b1010001: c <= 9'b1111100;
				8'b1010100: c <= 9'b1100110;
				8'b1100110: c <= 9'b100111;
				8'b101010: c <= 9'b100111001;
				8'b1011110: c <= 9'b110100001;
				8'b1100111: c <= 9'b111011110;
				8'b1011010: c <= 9'b110011001;
				8'b1000010: c <= 9'b110101010;
				8'b111101: c <= 9'b11101;
				8'b110000: c <= 9'b11011011;
				8'b111110: c <= 9'b1010101;
				8'b1100010: c <= 9'b110011101;
				8'b1110000: c <= 9'b111001111;
				8'b1101001: c <= 9'b100010001;
				8'b1110011: c <= 9'b101100010;
				8'b1001100: c <= 9'b1101111;
				8'b100001: c <= 9'b111110001;
				8'b1000110: c <= 9'b111000011;
				8'b1110010: c <= 9'b1001000;
				8'b1010000: c <= 9'b110001000;
				8'b1111010: c <= 9'b110011001;
				8'b1010101: c <= 9'b110110011;
				8'b111011: c <= 9'b100001001;
				8'b1001101: c <= 9'b10011111;
				8'b111111: c <= 9'b111011100;
				8'b1101110: c <= 9'b10010111;
				8'b1111011: c <= 9'b10110101;
				8'b1001011: c <= 9'b10101001;
				8'b1101111: c <= 9'b101001110;
				8'b1101000: c <= 9'b11011;
				8'b101100: c <= 9'b110111100;
				8'b100100: c <= 9'b101001111;
				8'b1111000: c <= 9'b100000101;
				8'b1000101: c <= 9'b1101110;
				8'b1011001: c <= 9'b111001011;
				8'b110100: c <= 9'b1011011;
				8'b1111001: c <= 9'b11100;
				8'b1110001: c <= 9'b11111000;
				8'b1001111: c <= 9'b10111000;
				8'b1100101: c <= 9'b110000011;
				8'b1111110: c <= 9'b111100001;
				8'b1111100: c <= 9'b1000111;
				8'b1010110: c <= 9'b101101101;
				8'b110010: c <= 9'b11000;
				8'b1101101: c <= 9'b111001010;
				8'b100011: c <= 9'b1010001;
				8'b1110101: c <= 9'b110011001;
				8'b1111101: c <= 9'b101001;
				8'b101001: c <= 9'b11;
				8'b1010010: c <= 9'b1100100;
				8'b1011000: c <= 9'b110000101;
				8'b101110: c <= 9'b10110;
				8'b1000001: c <= 9'b1110001;
				default: c <= 9'b0;
			endcase
			9'b100001101 : case(di)
				8'b1000011: c <= 9'b11101;
				8'b101000: c <= 9'b111101010;
				8'b111010: c <= 9'b110000110;
				8'b110110: c <= 9'b10001000;
				8'b1100100: c <= 9'b10110101;
				8'b1000000: c <= 9'b11001000;
				8'b1110110: c <= 9'b111010010;
				8'b100101: c <= 9'b110011100;
				8'b101111: c <= 9'b10111000;
				8'b100110: c <= 9'b11110011;
				8'b1100011: c <= 9'b111111001;
				8'b1001000: c <= 9'b101001001;
				8'b111000: c <= 9'b11001111;
				8'b110001: c <= 9'b101110110;
				8'b1010111: c <= 9'b111100101;
				8'b1001110: c <= 9'b10000110;
				8'b1101010: c <= 9'b110000101;
				8'b1001001: c <= 9'b1001110;
				8'b1100000: c <= 9'b100011100;
				8'b110111: c <= 9'b100110110;
				8'b1011101: c <= 9'b110000011;
				8'b1011011: c <= 9'b10101101;
				8'b111001: c <= 9'b11011100;
				8'b1001010: c <= 9'b101110101;
				8'b110011: c <= 9'b110001101;
				8'b1101100: c <= 9'b100010110;
				8'b1110111: c <= 9'b100000110;
				8'b101011: c <= 9'b10000110;
				8'b1101011: c <= 9'b11101000;
				8'b111100: c <= 9'b110110011;
				8'b1000111: c <= 9'b110011010;
				8'b1011111: c <= 9'b110100;
				8'b1110100: c <= 9'b101010110;
				8'b101101: c <= 9'b10110010;
				8'b1010011: c <= 9'b111110101;
				8'b1100001: c <= 9'b10000011;
				8'b110101: c <= 9'b11110111;
				8'b1000100: c <= 9'b1111000;
				8'b1010001: c <= 9'b10100010;
				8'b1010100: c <= 9'b101110010;
				8'b1100110: c <= 9'b10000011;
				8'b101010: c <= 9'b1010000;
				8'b1011110: c <= 9'b101011000;
				8'b1100111: c <= 9'b100000111;
				8'b1011010: c <= 9'b1;
				8'b1000010: c <= 9'b1100010;
				8'b111101: c <= 9'b111101000;
				8'b110000: c <= 9'b101001011;
				8'b111110: c <= 9'b100000001;
				8'b1100010: c <= 9'b100101111;
				8'b1110000: c <= 9'b100010100;
				8'b1101001: c <= 9'b110111111;
				8'b1110011: c <= 9'b11010100;
				8'b1001100: c <= 9'b11011001;
				8'b100001: c <= 9'b100100010;
				8'b1000110: c <= 9'b101100111;
				8'b1110010: c <= 9'b100011101;
				8'b1010000: c <= 9'b10111111;
				8'b1111010: c <= 9'b11110011;
				8'b1010101: c <= 9'b110000011;
				8'b111011: c <= 9'b1;
				8'b1001101: c <= 9'b1100;
				8'b111111: c <= 9'b110010001;
				8'b1101110: c <= 9'b110000111;
				8'b1111011: c <= 9'b101101101;
				8'b1001011: c <= 9'b111110000;
				8'b1101111: c <= 9'b10101100;
				8'b1101000: c <= 9'b110010101;
				8'b101100: c <= 9'b1000111;
				8'b100100: c <= 9'b10110101;
				8'b1111000: c <= 9'b100010110;
				8'b1000101: c <= 9'b10100100;
				8'b1011001: c <= 9'b11;
				8'b110100: c <= 9'b110011010;
				8'b1111001: c <= 9'b110111001;
				8'b1110001: c <= 9'b101000001;
				8'b1001111: c <= 9'b100110110;
				8'b1100101: c <= 9'b110001100;
				8'b1111110: c <= 9'b11111011;
				8'b1111100: c <= 9'b1001001;
				8'b1010110: c <= 9'b10000011;
				8'b110010: c <= 9'b101011010;
				8'b1101101: c <= 9'b100101111;
				8'b100011: c <= 9'b10111000;
				8'b1110101: c <= 9'b100100010;
				8'b1111101: c <= 9'b111010010;
				8'b101001: c <= 9'b10110011;
				8'b1010010: c <= 9'b111111111;
				8'b1011000: c <= 9'b11110;
				8'b101110: c <= 9'b100001100;
				8'b1000001: c <= 9'b1100001;
				default: c <= 9'b0;
			endcase
			9'b101010000 : case(di)
				8'b1000011: c <= 9'b110000110;
				8'b101000: c <= 9'b110100100;
				8'b111010: c <= 9'b1100101;
				8'b110110: c <= 9'b111110110;
				8'b1100100: c <= 9'b100100;
				8'b1000000: c <= 9'b110111111;
				8'b1110110: c <= 9'b100010110;
				8'b100101: c <= 9'b110011010;
				8'b101111: c <= 9'b11110100;
				8'b100110: c <= 9'b101011;
				8'b1100011: c <= 9'b100100011;
				8'b1001000: c <= 9'b111001;
				8'b111000: c <= 9'b10111001;
				8'b110001: c <= 9'b111000100;
				8'b1010111: c <= 9'b111011;
				8'b1001110: c <= 9'b110100101;
				8'b1101010: c <= 9'b101100;
				8'b1001001: c <= 9'b111011;
				8'b1100000: c <= 9'b100001101;
				8'b110111: c <= 9'b1011000;
				8'b1011101: c <= 9'b1100100;
				8'b1011011: c <= 9'b11011100;
				8'b111001: c <= 9'b110100001;
				8'b1001010: c <= 9'b111000000;
				8'b110011: c <= 9'b10;
				8'b1101100: c <= 9'b10100;
				8'b1110111: c <= 9'b1100100;
				8'b101011: c <= 9'b110011110;
				8'b1101011: c <= 9'b110011010;
				8'b111100: c <= 9'b1100010;
				8'b1000111: c <= 9'b101101001;
				8'b1011111: c <= 9'b110010001;
				8'b1110100: c <= 9'b101110011;
				8'b101101: c <= 9'b11101011;
				8'b1010011: c <= 9'b10010011;
				8'b1100001: c <= 9'b1011001;
				8'b110101: c <= 9'b101100111;
				8'b1000100: c <= 9'b10100;
				8'b1010001: c <= 9'b10110010;
				8'b1010100: c <= 9'b1010101;
				8'b1100110: c <= 9'b11110001;
				8'b101010: c <= 9'b111001;
				8'b1011110: c <= 9'b101100010;
				8'b1100111: c <= 9'b1100100;
				8'b1011010: c <= 9'b110001011;
				8'b1000010: c <= 9'b111000000;
				8'b111101: c <= 9'b101010101;
				8'b110000: c <= 9'b100110110;
				8'b111110: c <= 9'b110010001;
				8'b1100010: c <= 9'b111010001;
				8'b1110000: c <= 9'b1111110;
				8'b1101001: c <= 9'b1011100;
				8'b1110011: c <= 9'b101011010;
				8'b1001100: c <= 9'b110011100;
				8'b100001: c <= 9'b101010111;
				8'b1000110: c <= 9'b100010001;
				8'b1110010: c <= 9'b100011000;
				8'b1010000: c <= 9'b111110110;
				8'b1111010: c <= 9'b100100001;
				8'b1010101: c <= 9'b100000100;
				8'b111011: c <= 9'b11100000;
				8'b1001101: c <= 9'b1000000;
				8'b111111: c <= 9'b100111;
				8'b1101110: c <= 9'b100110011;
				8'b1111011: c <= 9'b10001101;
				8'b1001011: c <= 9'b101010;
				8'b1101111: c <= 9'b11110110;
				8'b1101000: c <= 9'b110111001;
				8'b101100: c <= 9'b100011000;
				8'b100100: c <= 9'b11110100;
				8'b1111000: c <= 9'b100101110;
				8'b1000101: c <= 9'b101110100;
				8'b1011001: c <= 9'b1110100;
				8'b110100: c <= 9'b1010010;
				8'b1111001: c <= 9'b11010;
				8'b1110001: c <= 9'b1000010;
				8'b1001111: c <= 9'b10000111;
				8'b1100101: c <= 9'b111101001;
				8'b1111110: c <= 9'b101000010;
				8'b1111100: c <= 9'b1011110;
				8'b1010110: c <= 9'b101001010;
				8'b110010: c <= 9'b10111000;
				8'b1101101: c <= 9'b11100011;
				8'b100011: c <= 9'b110100111;
				8'b1110101: c <= 9'b111010100;
				8'b1111101: c <= 9'b11101;
				8'b101001: c <= 9'b110101;
				8'b1010010: c <= 9'b100011100;
				8'b1011000: c <= 9'b111101100;
				8'b101110: c <= 9'b100000111;
				8'b1000001: c <= 9'b101101;
				default: c <= 9'b0;
			endcase
			9'b1111110 : case(di)
				8'b1000011: c <= 9'b11000;
				8'b101000: c <= 9'b10111011;
				8'b111010: c <= 9'b100;
				8'b110110: c <= 9'b10011000;
				8'b1100100: c <= 9'b10011111;
				8'b1000000: c <= 9'b101010;
				8'b1110110: c <= 9'b111100;
				8'b100101: c <= 9'b10011111;
				8'b101111: c <= 9'b10100111;
				8'b100110: c <= 9'b101010111;
				8'b1100011: c <= 9'b1011001;
				8'b1001000: c <= 9'b100001010;
				8'b111000: c <= 9'b11;
				8'b110001: c <= 9'b101000011;
				8'b1010111: c <= 9'b10110010;
				8'b1001110: c <= 9'b11100111;
				8'b1101010: c <= 9'b10110100;
				8'b1001001: c <= 9'b1000111;
				8'b1100000: c <= 9'b111010110;
				8'b110111: c <= 9'b101101110;
				8'b1011101: c <= 9'b100011;
				8'b1011011: c <= 9'b1001001;
				8'b111001: c <= 9'b101;
				8'b1001010: c <= 9'b110011111;
				8'b110011: c <= 9'b110011;
				8'b1101100: c <= 9'b100011001;
				8'b1110111: c <= 9'b1011100;
				8'b101011: c <= 9'b101010010;
				8'b1101011: c <= 9'b111001010;
				8'b111100: c <= 9'b110000000;
				8'b1000111: c <= 9'b100010;
				8'b1011111: c <= 9'b10110110;
				8'b1110100: c <= 9'b111011101;
				8'b101101: c <= 9'b100110101;
				8'b1010011: c <= 9'b11111100;
				8'b1100001: c <= 9'b1111010;
				8'b110101: c <= 9'b101110010;
				8'b1000100: c <= 9'b100100101;
				8'b1010001: c <= 9'b11000011;
				8'b1010100: c <= 9'b11011;
				8'b1100110: c <= 9'b110101111;
				8'b101010: c <= 9'b1111111;
				8'b1011110: c <= 9'b1111;
				8'b1100111: c <= 9'b111111101;
				8'b1011010: c <= 9'b101100101;
				8'b1000010: c <= 9'b101110010;
				8'b111101: c <= 9'b10001101;
				8'b110000: c <= 9'b110100;
				8'b111110: c <= 9'b1110011;
				8'b1100010: c <= 9'b101010001;
				8'b1110000: c <= 9'b110110100;
				8'b1101001: c <= 9'b110001011;
				8'b1110011: c <= 9'b11111;
				8'b1001100: c <= 9'b10001010;
				8'b100001: c <= 9'b110001000;
				8'b1000110: c <= 9'b1110001;
				8'b1110010: c <= 9'b11011110;
				8'b1010000: c <= 9'b100110011;
				8'b1111010: c <= 9'b100111;
				8'b1010101: c <= 9'b1101100;
				8'b111011: c <= 9'b101110000;
				8'b1001101: c <= 9'b11001110;
				8'b111111: c <= 9'b111000;
				8'b1101110: c <= 9'b1110111;
				8'b1111011: c <= 9'b101000011;
				8'b1001011: c <= 9'b11111100;
				8'b1101111: c <= 9'b1101110;
				8'b1101000: c <= 9'b10010101;
				8'b101100: c <= 9'b1110010;
				8'b100100: c <= 9'b10010;
				8'b1111000: c <= 9'b111100011;
				8'b1000101: c <= 9'b101110110;
				8'b1011001: c <= 9'b110011000;
				8'b110100: c <= 9'b110010100;
				8'b1111001: c <= 9'b110011111;
				8'b1110001: c <= 9'b10100011;
				8'b1001111: c <= 9'b11001;
				8'b1100101: c <= 9'b111101001;
				8'b1111110: c <= 9'b11101101;
				8'b1111100: c <= 9'b101010101;
				8'b1010110: c <= 9'b110100110;
				8'b110010: c <= 9'b100110110;
				8'b1101101: c <= 9'b110010110;
				8'b100011: c <= 9'b100001011;
				8'b1110101: c <= 9'b11111000;
				8'b1111101: c <= 9'b110001001;
				8'b101001: c <= 9'b11111101;
				8'b1010010: c <= 9'b100011001;
				8'b1011000: c <= 9'b111110011;
				8'b101110: c <= 9'b100101001;
				8'b1000001: c <= 9'b100011001;
				default: c <= 9'b0;
			endcase
			9'b10010 : case(di)
				8'b1000011: c <= 9'b11000010;
				8'b101000: c <= 9'b11110101;
				8'b111010: c <= 9'b101010111;
				8'b110110: c <= 9'b1100110;
				8'b1100100: c <= 9'b11111101;
				8'b1000000: c <= 9'b100010110;
				8'b1110110: c <= 9'b11;
				8'b100101: c <= 9'b101101100;
				8'b101111: c <= 9'b100110110;
				8'b100110: c <= 9'b1000100;
				8'b1100011: c <= 9'b100110100;
				8'b1001000: c <= 9'b10010100;
				8'b111000: c <= 9'b100000110;
				8'b110001: c <= 9'b100101010;
				8'b1010111: c <= 9'b101010001;
				8'b1001110: c <= 9'b1111111;
				8'b1101010: c <= 9'b111010000;
				8'b1001001: c <= 9'b11110110;
				8'b1100000: c <= 9'b111110000;
				8'b110111: c <= 9'b11000011;
				8'b1011101: c <= 9'b100011011;
				8'b1011011: c <= 9'b11010001;
				8'b111001: c <= 9'b1010110;
				8'b1001010: c <= 9'b111110000;
				8'b110011: c <= 9'b1111101;
				8'b1101100: c <= 9'b100111110;
				8'b1110111: c <= 9'b111110110;
				8'b101011: c <= 9'b101001;
				8'b1101011: c <= 9'b11110110;
				8'b111100: c <= 9'b100010000;
				8'b1000111: c <= 9'b100110000;
				8'b1011111: c <= 9'b110011110;
				8'b1110100: c <= 9'b101111000;
				8'b101101: c <= 9'b101110;
				8'b1010011: c <= 9'b111;
				8'b1100001: c <= 9'b10111011;
				8'b110101: c <= 9'b11001101;
				8'b1000100: c <= 9'b1000111;
				8'b1010001: c <= 9'b111111011;
				8'b1010100: c <= 9'b1110101;
				8'b1100110: c <= 9'b111100;
				8'b101010: c <= 9'b10010;
				8'b1011110: c <= 9'b111011110;
				8'b1100111: c <= 9'b101011110;
				8'b1011010: c <= 9'b10001110;
				8'b1000010: c <= 9'b1101001;
				8'b111101: c <= 9'b111011001;
				8'b110000: c <= 9'b1110101;
				8'b111110: c <= 9'b100100001;
				8'b1100010: c <= 9'b100101000;
				8'b1110000: c <= 9'b111100100;
				8'b1101001: c <= 9'b110101001;
				8'b1110011: c <= 9'b100100101;
				8'b1001100: c <= 9'b11101100;
				8'b100001: c <= 9'b1000110;
				8'b1000110: c <= 9'b10011101;
				8'b1110010: c <= 9'b100101;
				8'b1010000: c <= 9'b101010011;
				8'b1111010: c <= 9'b100010011;
				8'b1010101: c <= 9'b10011100;
				8'b111011: c <= 9'b110101001;
				8'b1001101: c <= 9'b110011101;
				8'b111111: c <= 9'b11001101;
				8'b1101110: c <= 9'b11000;
				8'b1111011: c <= 9'b10001101;
				8'b1001011: c <= 9'b111000101;
				8'b1101111: c <= 9'b10100101;
				8'b1101000: c <= 9'b10011;
				8'b101100: c <= 9'b110111100;
				8'b100100: c <= 9'b110110111;
				8'b1111000: c <= 9'b101100001;
				8'b1000101: c <= 9'b111000010;
				8'b1011001: c <= 9'b110000010;
				8'b110100: c <= 9'b101010111;
				8'b1111001: c <= 9'b101001011;
				8'b1110001: c <= 9'b1111011;
				8'b1001111: c <= 9'b111101000;
				8'b1100101: c <= 9'b101001010;
				8'b1111110: c <= 9'b100110111;
				8'b1111100: c <= 9'b110100010;
				8'b1010110: c <= 9'b110111110;
				8'b110010: c <= 9'b111111000;
				8'b1101101: c <= 9'b110000111;
				8'b100011: c <= 9'b10010000;
				8'b1110101: c <= 9'b111001101;
				8'b1111101: c <= 9'b101111010;
				8'b101001: c <= 9'b110100111;
				8'b1010010: c <= 9'b101001010;
				8'b1011000: c <= 9'b10100111;
				8'b101110: c <= 9'b101101101;
				8'b1000001: c <= 9'b101101010;
				default: c <= 9'b0;
			endcase
			9'b111011100 : case(di)
				8'b1000011: c <= 9'b100010;
				8'b101000: c <= 9'b10111001;
				8'b111010: c <= 9'b101100010;
				8'b110110: c <= 9'b10010001;
				8'b1100100: c <= 9'b111011111;
				8'b1000000: c <= 9'b110011000;
				8'b1110110: c <= 9'b100010110;
				8'b100101: c <= 9'b100010110;
				8'b101111: c <= 9'b100101110;
				8'b100110: c <= 9'b111010001;
				8'b1100011: c <= 9'b100011001;
				8'b1001000: c <= 9'b11110000;
				8'b111000: c <= 9'b110101110;
				8'b110001: c <= 9'b110011;
				8'b1010111: c <= 9'b11001111;
				8'b1001110: c <= 9'b10111;
				8'b1101010: c <= 9'b100101101;
				8'b1001001: c <= 9'b11101011;
				8'b1100000: c <= 9'b101101011;
				8'b110111: c <= 9'b110111111;
				8'b1011101: c <= 9'b1010110;
				8'b1011011: c <= 9'b110011010;
				8'b111001: c <= 9'b110101101;
				8'b1001010: c <= 9'b110111011;
				8'b110011: c <= 9'b111111;
				8'b1101100: c <= 9'b101110110;
				8'b1110111: c <= 9'b1111010;
				8'b101011: c <= 9'b1110101;
				8'b1101011: c <= 9'b100011000;
				8'b111100: c <= 9'b100;
				8'b1000111: c <= 9'b11100001;
				8'b1011111: c <= 9'b10101010;
				8'b1110100: c <= 9'b11011110;
				8'b101101: c <= 9'b101101001;
				8'b1010011: c <= 9'b1001011;
				8'b1100001: c <= 9'b111011;
				8'b110101: c <= 9'b110001111;
				8'b1000100: c <= 9'b1100101;
				8'b1010001: c <= 9'b11001101;
				8'b1010100: c <= 9'b1110101;
				8'b1100110: c <= 9'b1110000;
				8'b101010: c <= 9'b10001100;
				8'b1011110: c <= 9'b100001111;
				8'b1100111: c <= 9'b100101100;
				8'b1011010: c <= 9'b1100110;
				8'b1000010: c <= 9'b10111101;
				8'b111101: c <= 9'b111010010;
				8'b110000: c <= 9'b1110;
				8'b111110: c <= 9'b101100000;
				8'b1100010: c <= 9'b100101110;
				8'b1110000: c <= 9'b110010;
				8'b1101001: c <= 9'b101100100;
				8'b1110011: c <= 9'b100011101;
				8'b1001100: c <= 9'b1111;
				8'b100001: c <= 9'b111000011;
				8'b1000110: c <= 9'b110111011;
				8'b1110010: c <= 9'b110000011;
				8'b1010000: c <= 9'b100110110;
				8'b1111010: c <= 9'b10000111;
				8'b1010101: c <= 9'b10101101;
				8'b111011: c <= 9'b100111110;
				8'b1001101: c <= 9'b1001100;
				8'b111111: c <= 9'b10101101;
				8'b1101110: c <= 9'b111110110;
				8'b1111011: c <= 9'b110111010;
				8'b1001011: c <= 9'b11010001;
				8'b1101111: c <= 9'b100011011;
				8'b1101000: c <= 9'b111011100;
				8'b101100: c <= 9'b10110001;
				8'b100100: c <= 9'b11000011;
				8'b1111000: c <= 9'b111111111;
				8'b1000101: c <= 9'b111001101;
				8'b1011001: c <= 9'b10110;
				8'b110100: c <= 9'b10101100;
				8'b1111001: c <= 9'b100010011;
				8'b1110001: c <= 9'b11101;
				8'b1001111: c <= 9'b111101010;
				8'b1100101: c <= 9'b111111110;
				8'b1111110: c <= 9'b101101000;
				8'b1111100: c <= 9'b1100000;
				8'b1010110: c <= 9'b10101011;
				8'b110010: c <= 9'b110011111;
				8'b1101101: c <= 9'b101101110;
				8'b100011: c <= 9'b101110001;
				8'b1110101: c <= 9'b110111001;
				8'b1111101: c <= 9'b10111111;
				8'b101001: c <= 9'b100111010;
				8'b1010010: c <= 9'b10110010;
				8'b1011000: c <= 9'b10110010;
				8'b101110: c <= 9'b1100010;
				8'b1000001: c <= 9'b10010111;
				default: c <= 9'b0;
			endcase
			9'b100110010 : case(di)
				8'b1000011: c <= 9'b110011011;
				8'b101000: c <= 9'b1111;
				8'b111010: c <= 9'b110110110;
				8'b110110: c <= 9'b111101101;
				8'b1100100: c <= 9'b111010110;
				8'b1000000: c <= 9'b11101001;
				8'b1110110: c <= 9'b1111110;
				8'b100101: c <= 9'b10000110;
				8'b101111: c <= 9'b10000000;
				8'b100110: c <= 9'b10111111;
				8'b1100011: c <= 9'b11010100;
				8'b1001000: c <= 9'b100111111;
				8'b111000: c <= 9'b110001;
				8'b110001: c <= 9'b10011010;
				8'b1010111: c <= 9'b1111;
				8'b1001110: c <= 9'b1010000;
				8'b1101010: c <= 9'b1101101;
				8'b1001001: c <= 9'b11010001;
				8'b1100000: c <= 9'b111000101;
				8'b110111: c <= 9'b11100011;
				8'b1011101: c <= 9'b110100010;
				8'b1011011: c <= 9'b101110011;
				8'b111001: c <= 9'b11011101;
				8'b1001010: c <= 9'b10000110;
				8'b110011: c <= 9'b1110;
				8'b1101100: c <= 9'b10000010;
				8'b1110111: c <= 9'b11101101;
				8'b101011: c <= 9'b101111000;
				8'b1101011: c <= 9'b10111110;
				8'b111100: c <= 9'b111000100;
				8'b1000111: c <= 9'b100111010;
				8'b1011111: c <= 9'b111100111;
				8'b1110100: c <= 9'b110101011;
				8'b101101: c <= 9'b10000000;
				8'b1010011: c <= 9'b111010100;
				8'b1100001: c <= 9'b11010010;
				8'b110101: c <= 9'b100010100;
				8'b1000100: c <= 9'b1111101;
				8'b1010001: c <= 9'b11011011;
				8'b1010100: c <= 9'b101000;
				8'b1100110: c <= 9'b110000010;
				8'b101010: c <= 9'b10100000;
				8'b1011110: c <= 9'b100101111;
				8'b1100111: c <= 9'b100111;
				8'b1011010: c <= 9'b11010111;
				8'b1000010: c <= 9'b1111101;
				8'b111101: c <= 9'b11101100;
				8'b110000: c <= 9'b101010011;
				8'b111110: c <= 9'b10001100;
				8'b1100010: c <= 9'b100111011;
				8'b1110000: c <= 9'b1100010;
				8'b1101001: c <= 9'b111010000;
				8'b1110011: c <= 9'b110100;
				8'b1001100: c <= 9'b10000011;
				8'b100001: c <= 9'b110101;
				8'b1000110: c <= 9'b10010100;
				8'b1110010: c <= 9'b1010010;
				8'b1010000: c <= 9'b10110110;
				8'b1111010: c <= 9'b1111101;
				8'b1010101: c <= 9'b1000011;
				8'b111011: c <= 9'b110010010;
				8'b1001101: c <= 9'b100001011;
				8'b111111: c <= 9'b111111101;
				8'b1101110: c <= 9'b111110011;
				8'b1111011: c <= 9'b1110101;
				8'b1001011: c <= 9'b110101;
				8'b1101111: c <= 9'b11011110;
				8'b1101000: c <= 9'b100111010;
				8'b101100: c <= 9'b100111010;
				8'b100100: c <= 9'b1101101;
				8'b1111000: c <= 9'b11110;
				8'b1000101: c <= 9'b110000000;
				8'b1011001: c <= 9'b111001011;
				8'b110100: c <= 9'b110111110;
				8'b1111001: c <= 9'b101010000;
				8'b1110001: c <= 9'b1100001;
				8'b1001111: c <= 9'b110110101;
				8'b1100101: c <= 9'b111011100;
				8'b1111110: c <= 9'b10011;
				8'b1111100: c <= 9'b1101110;
				8'b1010110: c <= 9'b101011000;
				8'b110010: c <= 9'b11010100;
				8'b1101101: c <= 9'b101001111;
				8'b100011: c <= 9'b111010110;
				8'b1110101: c <= 9'b111011100;
				8'b1111101: c <= 9'b101101011;
				8'b101001: c <= 9'b100011001;
				8'b1010010: c <= 9'b101100110;
				8'b1011000: c <= 9'b110000101;
				8'b101110: c <= 9'b100101110;
				8'b1000001: c <= 9'b100010011;
				default: c <= 9'b0;
			endcase
			9'b101000011 : case(di)
				8'b1000011: c <= 9'b101110101;
				8'b101000: c <= 9'b11001000;
				8'b111010: c <= 9'b10001010;
				8'b110110: c <= 9'b100010011;
				8'b1100100: c <= 9'b101010011;
				8'b1000000: c <= 9'b101001011;
				8'b1110110: c <= 9'b10000110;
				8'b100101: c <= 9'b10100101;
				8'b101111: c <= 9'b1001010;
				8'b100110: c <= 9'b111010100;
				8'b1100011: c <= 9'b10011;
				8'b1001000: c <= 9'b11100101;
				8'b111000: c <= 9'b1101001;
				8'b110001: c <= 9'b110010001;
				8'b1010111: c <= 9'b10101110;
				8'b1001110: c <= 9'b110011100;
				8'b1101010: c <= 9'b111100101;
				8'b1001001: c <= 9'b1011111;
				8'b1100000: c <= 9'b11001110;
				8'b110111: c <= 9'b10100111;
				8'b1011101: c <= 9'b10001111;
				8'b1011011: c <= 9'b1111111;
				8'b111001: c <= 9'b1111011;
				8'b1001010: c <= 9'b111100001;
				8'b110011: c <= 9'b111111110;
				8'b1101100: c <= 9'b111100011;
				8'b1110111: c <= 9'b1010111;
				8'b101011: c <= 9'b111110110;
				8'b1101011: c <= 9'b111101111;
				8'b111100: c <= 9'b10101111;
				8'b1000111: c <= 9'b10110011;
				8'b1011111: c <= 9'b1010101;
				8'b1110100: c <= 9'b101001001;
				8'b101101: c <= 9'b1011011;
				8'b1010011: c <= 9'b100110;
				8'b1100001: c <= 9'b1011110;
				8'b110101: c <= 9'b10011001;
				8'b1000100: c <= 9'b110000101;
				8'b1010001: c <= 9'b1101000;
				8'b1010100: c <= 9'b110111001;
				8'b1100110: c <= 9'b110011010;
				8'b101010: c <= 9'b1010101;
				8'b1011110: c <= 9'b101111111;
				8'b1100111: c <= 9'b101;
				8'b1011010: c <= 9'b1000100;
				8'b1000010: c <= 9'b110111011;
				8'b111101: c <= 9'b100001;
				8'b110000: c <= 9'b110001010;
				8'b111110: c <= 9'b10111111;
				8'b1100010: c <= 9'b101010000;
				8'b1110000: c <= 9'b10010;
				8'b1101001: c <= 9'b101110110;
				8'b1110011: c <= 9'b100101010;
				8'b1001100: c <= 9'b10010111;
				8'b100001: c <= 9'b1001100;
				8'b1000110: c <= 9'b1111100;
				8'b1110010: c <= 9'b10011011;
				8'b1010000: c <= 9'b10110001;
				8'b1111010: c <= 9'b10010011;
				8'b1010101: c <= 9'b100000001;
				8'b111011: c <= 9'b111001101;
				8'b1001101: c <= 9'b110011010;
				8'b111111: c <= 9'b1100011;
				8'b1101110: c <= 9'b110010010;
				8'b1111011: c <= 9'b101101010;
				8'b1001011: c <= 9'b110100100;
				8'b1101111: c <= 9'b11110001;
				8'b1101000: c <= 9'b100011001;
				8'b101100: c <= 9'b1100110;
				8'b100100: c <= 9'b111001110;
				8'b1111000: c <= 9'b10100000;
				8'b1000101: c <= 9'b1101111;
				8'b1011001: c <= 9'b10001101;
				8'b110100: c <= 9'b11011101;
				8'b1111001: c <= 9'b111011010;
				8'b1110001: c <= 9'b111000110;
				8'b1001111: c <= 9'b100111;
				8'b1100101: c <= 9'b11101100;
				8'b1111110: c <= 9'b110000110;
				8'b1111100: c <= 9'b110101100;
				8'b1010110: c <= 9'b110000;
				8'b110010: c <= 9'b101111001;
				8'b1101101: c <= 9'b10101001;
				8'b100011: c <= 9'b100000110;
				8'b1110101: c <= 9'b10101;
				8'b1111101: c <= 9'b10001011;
				8'b101001: c <= 9'b111100011;
				8'b1010010: c <= 9'b101011010;
				8'b1011000: c <= 9'b101110101;
				8'b101110: c <= 9'b1111011;
				8'b1000001: c <= 9'b101100011;
				default: c <= 9'b0;
			endcase
			9'b111 : case(di)
				8'b1000011: c <= 9'b10111010;
				8'b101000: c <= 9'b1011100;
				8'b111010: c <= 9'b100110010;
				8'b110110: c <= 9'b111010111;
				8'b1100100: c <= 9'b110001011;
				8'b1000000: c <= 9'b111011010;
				8'b1110110: c <= 9'b100011101;
				8'b100101: c <= 9'b101110011;
				8'b101111: c <= 9'b100000011;
				8'b100110: c <= 9'b1111001;
				8'b1100011: c <= 9'b100010111;
				8'b1001000: c <= 9'b110000110;
				8'b111000: c <= 9'b100001001;
				8'b110001: c <= 9'b110011000;
				8'b1010111: c <= 9'b1000010;
				8'b1001110: c <= 9'b111101101;
				8'b1101010: c <= 9'b110110100;
				8'b1001001: c <= 9'b101011;
				8'b1100000: c <= 9'b101101011;
				8'b110111: c <= 9'b100011001;
				8'b1011101: c <= 9'b111000011;
				8'b1011011: c <= 9'b11100101;
				8'b111001: c <= 9'b1100010;
				8'b1001010: c <= 9'b1;
				8'b110011: c <= 9'b111000101;
				8'b1101100: c <= 9'b1010000;
				8'b1110111: c <= 9'b10001111;
				8'b101011: c <= 9'b101011000;
				8'b1101011: c <= 9'b11001011;
				8'b111100: c <= 9'b11001010;
				8'b1000111: c <= 9'b1111;
				8'b1011111: c <= 9'b100000010;
				8'b1110100: c <= 9'b11011000;
				8'b101101: c <= 9'b10111010;
				8'b1010011: c <= 9'b111101010;
				8'b1100001: c <= 9'b110100101;
				8'b110101: c <= 9'b111110001;
				8'b1000100: c <= 9'b11110101;
				8'b1010001: c <= 9'b111111111;
				8'b1010100: c <= 9'b10100111;
				8'b1100110: c <= 9'b11110010;
				8'b101010: c <= 9'b110010001;
				8'b1011110: c <= 9'b100110110;
				8'b1100111: c <= 9'b11101001;
				8'b1011010: c <= 9'b110110010;
				8'b1000010: c <= 9'b11100;
				8'b111101: c <= 9'b101100;
				8'b110000: c <= 9'b1001011;
				8'b111110: c <= 9'b101010100;
				8'b1100010: c <= 9'b1101100;
				8'b1110000: c <= 9'b110001100;
				8'b1101001: c <= 9'b10101101;
				8'b1110011: c <= 9'b101101001;
				8'b1001100: c <= 9'b101101011;
				8'b100001: c <= 9'b1111000;
				8'b1000110: c <= 9'b11000111;
				8'b1110010: c <= 9'b11110101;
				8'b1010000: c <= 9'b11000100;
				8'b1111010: c <= 9'b1110000;
				8'b1010101: c <= 9'b110000111;
				8'b111011: c <= 9'b101011110;
				8'b1001101: c <= 9'b100101001;
				8'b111111: c <= 9'b110000;
				8'b1101110: c <= 9'b1111010;
				8'b1111011: c <= 9'b101110001;
				8'b1001011: c <= 9'b110100011;
				8'b1101111: c <= 9'b100110010;
				8'b1101000: c <= 9'b100111010;
				8'b101100: c <= 9'b1011010;
				8'b100100: c <= 9'b111010000;
				8'b1111000: c <= 9'b111100010;
				8'b1000101: c <= 9'b10000101;
				8'b1011001: c <= 9'b100111010;
				8'b110100: c <= 9'b10000101;
				8'b1111001: c <= 9'b100110;
				8'b1110001: c <= 9'b111011100;
				8'b1001111: c <= 9'b100011;
				8'b1100101: c <= 9'b1111100;
				8'b1111110: c <= 9'b100101110;
				8'b1111100: c <= 9'b11000001;
				8'b1010110: c <= 9'b10100;
				8'b110010: c <= 9'b111001;
				8'b1101101: c <= 9'b100011111;
				8'b100011: c <= 9'b111010111;
				8'b1110101: c <= 9'b111001101;
				8'b1111101: c <= 9'b111001;
				8'b101001: c <= 9'b1111101;
				8'b1010010: c <= 9'b11010101;
				8'b1011000: c <= 9'b10011001;
				8'b101110: c <= 9'b110101010;
				8'b1000001: c <= 9'b101110111;
				default: c <= 9'b0;
			endcase
			9'b1100000 : case(di)
				8'b1000011: c <= 9'b111111000;
				8'b101000: c <= 9'b11000111;
				8'b111010: c <= 9'b11000110;
				8'b110110: c <= 9'b11000011;
				8'b1100100: c <= 9'b10001000;
				8'b1000000: c <= 9'b101100001;
				8'b1110110: c <= 9'b100001100;
				8'b100101: c <= 9'b111011010;
				8'b101111: c <= 9'b1111110;
				8'b100110: c <= 9'b110101110;
				8'b1100011: c <= 9'b101011001;
				8'b1001000: c <= 9'b11;
				8'b111000: c <= 9'b1111001;
				8'b110001: c <= 9'b110101;
				8'b1010111: c <= 9'b110010010;
				8'b1001110: c <= 9'b10;
				8'b1101010: c <= 9'b1011001;
				8'b1001001: c <= 9'b11;
				8'b1100000: c <= 9'b101001011;
				8'b110111: c <= 9'b111100000;
				8'b1011101: c <= 9'b11010001;
				8'b1011011: c <= 9'b110101100;
				8'b111001: c <= 9'b110100111;
				8'b1001010: c <= 9'b1111101;
				8'b110011: c <= 9'b1001101;
				8'b1101100: c <= 9'b1011;
				8'b1110111: c <= 9'b100101010;
				8'b101011: c <= 9'b10001001;
				8'b1101011: c <= 9'b11000000;
				8'b111100: c <= 9'b10011011;
				8'b1000111: c <= 9'b1001001;
				8'b1011111: c <= 9'b111011001;
				8'b1110100: c <= 9'b110000;
				8'b101101: c <= 9'b111;
				8'b1010011: c <= 9'b100011100;
				8'b1100001: c <= 9'b101011001;
				8'b110101: c <= 9'b111111000;
				8'b1000100: c <= 9'b10000010;
				8'b1010001: c <= 9'b11100010;
				8'b1010100: c <= 9'b1111011;
				8'b1100110: c <= 9'b101;
				8'b101010: c <= 9'b1101100;
				8'b1011110: c <= 9'b11010001;
				8'b1100111: c <= 9'b101011110;
				8'b1011010: c <= 9'b1101000;
				8'b1000010: c <= 9'b111111101;
				8'b111101: c <= 9'b1110010;
				8'b110000: c <= 9'b110110010;
				8'b111110: c <= 9'b10010;
				8'b1100010: c <= 9'b110100000;
				8'b1110000: c <= 9'b100001111;
				8'b1101001: c <= 9'b100011111;
				8'b1110011: c <= 9'b101001010;
				8'b1001100: c <= 9'b1001001;
				8'b100001: c <= 9'b101000;
				8'b1000110: c <= 9'b110011011;
				8'b1110010: c <= 9'b1101110;
				8'b1010000: c <= 9'b1100010;
				8'b1111010: c <= 9'b110010101;
				8'b1010101: c <= 9'b100001;
				8'b111011: c <= 9'b101010000;
				8'b1001101: c <= 9'b10000110;
				8'b111111: c <= 9'b11000001;
				8'b1101110: c <= 9'b111111010;
				8'b1111011: c <= 9'b1101110;
				8'b1001011: c <= 9'b10000110;
				8'b1101111: c <= 9'b100110100;
				8'b1101000: c <= 9'b101010;
				8'b101100: c <= 9'b111111001;
				8'b100100: c <= 9'b100101111;
				8'b1111000: c <= 9'b1010001;
				8'b1000101: c <= 9'b11000111;
				8'b1011001: c <= 9'b10111100;
				8'b110100: c <= 9'b110011111;
				8'b1111001: c <= 9'b111111010;
				8'b1110001: c <= 9'b100110;
				8'b1001111: c <= 9'b11101101;
				8'b1100101: c <= 9'b100101010;
				8'b1111110: c <= 9'b110001001;
				8'b1111100: c <= 9'b100100010;
				8'b1010110: c <= 9'b1111001;
				8'b110010: c <= 9'b101110111;
				8'b1101101: c <= 9'b11000100;
				8'b100011: c <= 9'b110100;
				8'b1110101: c <= 9'b111100;
				8'b1111101: c <= 9'b111100110;
				8'b101001: c <= 9'b1010000;
				8'b1010010: c <= 9'b110101;
				8'b1011000: c <= 9'b10100101;
				8'b101110: c <= 9'b101111110;
				8'b1000001: c <= 9'b101111001;
				default: c <= 9'b0;
			endcase
			9'b1100110 : case(di)
				8'b1000011: c <= 9'b10111001;
				8'b101000: c <= 9'b111101101;
				8'b111010: c <= 9'b11010101;
				8'b110110: c <= 9'b100010000;
				8'b1100100: c <= 9'b101101011;
				8'b1000000: c <= 9'b10101101;
				8'b1110110: c <= 9'b110011110;
				8'b100101: c <= 9'b110011111;
				8'b101111: c <= 9'b10100111;
				8'b100110: c <= 9'b1111001;
				8'b1100011: c <= 9'b1100011;
				8'b1001000: c <= 9'b11001110;
				8'b111000: c <= 9'b111001111;
				8'b110001: c <= 9'b10011101;
				8'b1010111: c <= 9'b11001000;
				8'b1001110: c <= 9'b111001000;
				8'b1101010: c <= 9'b101110100;
				8'b1001001: c <= 9'b111101001;
				8'b1100000: c <= 9'b11001010;
				8'b110111: c <= 9'b1000000;
				8'b1011101: c <= 9'b10101111;
				8'b1011011: c <= 9'b11000111;
				8'b111001: c <= 9'b110000001;
				8'b1001010: c <= 9'b111101001;
				8'b110011: c <= 9'b11011;
				8'b1101100: c <= 9'b1100011;
				8'b1110111: c <= 9'b11011011;
				8'b101011: c <= 9'b1000100;
				8'b1101011: c <= 9'b101110011;
				8'b111100: c <= 9'b11010001;
				8'b1000111: c <= 9'b10110;
				8'b1011111: c <= 9'b101111000;
				8'b1110100: c <= 9'b110100;
				8'b101101: c <= 9'b110110;
				8'b1010011: c <= 9'b111000111;
				8'b1100001: c <= 9'b10011101;
				8'b110101: c <= 9'b11001101;
				8'b1000100: c <= 9'b10101010;
				8'b1010001: c <= 9'b111110001;
				8'b1010100: c <= 9'b110111010;
				8'b1100110: c <= 9'b11011101;
				8'b101010: c <= 9'b11001011;
				8'b1011110: c <= 9'b11100110;
				8'b1100111: c <= 9'b100101001;
				8'b1011010: c <= 9'b10101101;
				8'b1000010: c <= 9'b111111001;
				8'b111101: c <= 9'b101111001;
				8'b110000: c <= 9'b1111101;
				8'b111110: c <= 9'b100010100;
				8'b1100010: c <= 9'b1101000;
				8'b1110000: c <= 9'b10010;
				8'b1101001: c <= 9'b11001011;
				8'b1110011: c <= 9'b1011110;
				8'b1001100: c <= 9'b100110100;
				8'b100001: c <= 9'b111011011;
				8'b1000110: c <= 9'b10010000;
				8'b1110010: c <= 9'b11101011;
				8'b1010000: c <= 9'b10011101;
				8'b1111010: c <= 9'b100000000;
				8'b1010101: c <= 9'b11011110;
				8'b111011: c <= 9'b11001;
				8'b1001101: c <= 9'b100011010;
				8'b111111: c <= 9'b11000110;
				8'b1101110: c <= 9'b10100011;
				8'b1111011: c <= 9'b1110010;
				8'b1001011: c <= 9'b100110110;
				8'b1101111: c <= 9'b110100100;
				8'b1101000: c <= 9'b1001000;
				8'b101100: c <= 9'b10000101;
				8'b100100: c <= 9'b101111111;
				8'b1111000: c <= 9'b111100000;
				8'b1000101: c <= 9'b11011;
				8'b1011001: c <= 9'b10000110;
				8'b110100: c <= 9'b11000110;
				8'b1111001: c <= 9'b100110011;
				8'b1110001: c <= 9'b10010110;
				8'b1001111: c <= 9'b11011100;
				8'b1100101: c <= 9'b101100101;
				8'b1111110: c <= 9'b100010;
				8'b1111100: c <= 9'b11101111;
				8'b1010110: c <= 9'b100000011;
				8'b110010: c <= 9'b11001001;
				8'b1101101: c <= 9'b11101111;
				8'b100011: c <= 9'b10100101;
				8'b1110101: c <= 9'b1010000;
				8'b1111101: c <= 9'b101010010;
				8'b101001: c <= 9'b111001000;
				8'b1010010: c <= 9'b101010101;
				8'b1011000: c <= 9'b110000110;
				8'b101110: c <= 9'b101110100;
				8'b1000001: c <= 9'b1001;
				default: c <= 9'b0;
			endcase
			9'b11000100 : case(di)
				8'b1000011: c <= 9'b100010100;
				8'b101000: c <= 9'b1110;
				8'b111010: c <= 9'b100101011;
				8'b110110: c <= 9'b110100000;
				8'b1100100: c <= 9'b111011010;
				8'b1000000: c <= 9'b1;
				8'b1110110: c <= 9'b110000011;
				8'b100101: c <= 9'b111000;
				8'b101111: c <= 9'b101101110;
				8'b100110: c <= 9'b101101;
				8'b1100011: c <= 9'b1101010;
				8'b1001000: c <= 9'b111100100;
				8'b111000: c <= 9'b100111000;
				8'b110001: c <= 9'b1110;
				8'b1010111: c <= 9'b10101001;
				8'b1001110: c <= 9'b10010110;
				8'b1101010: c <= 9'b11100011;
				8'b1001001: c <= 9'b100101011;
				8'b1100000: c <= 9'b111011100;
				8'b110111: c <= 9'b1011100;
				8'b1011101: c <= 9'b101010;
				8'b1011011: c <= 9'b110111011;
				8'b111001: c <= 9'b110101100;
				8'b1001010: c <= 9'b11110001;
				8'b110011: c <= 9'b11000100;
				8'b1101100: c <= 9'b11111011;
				8'b1110111: c <= 9'b10110100;
				8'b101011: c <= 9'b1010011;
				8'b1101011: c <= 9'b110100;
				8'b111100: c <= 9'b11000011;
				8'b1000111: c <= 9'b10010;
				8'b1011111: c <= 9'b10010110;
				8'b1110100: c <= 9'b10110;
				8'b101101: c <= 9'b10011011;
				8'b1010011: c <= 9'b1001101;
				8'b1100001: c <= 9'b1111101;
				8'b110101: c <= 9'b101100;
				8'b1000100: c <= 9'b1101100;
				8'b1010001: c <= 9'b10000;
				8'b1010100: c <= 9'b111111010;
				8'b1100110: c <= 9'b11101011;
				8'b101010: c <= 9'b100000010;
				8'b1011110: c <= 9'b1111011;
				8'b1100111: c <= 9'b1110;
				8'b1011010: c <= 9'b110001100;
				8'b1000010: c <= 9'b10011000;
				8'b111101: c <= 9'b1101110;
				8'b110000: c <= 9'b10101011;
				8'b111110: c <= 9'b1110111;
				8'b1100010: c <= 9'b111101000;
				8'b1110000: c <= 9'b110001111;
				8'b1101001: c <= 9'b111101110;
				8'b1110011: c <= 9'b110110010;
				8'b1001100: c <= 9'b110100011;
				8'b100001: c <= 9'b100111111;
				8'b1000110: c <= 9'b10001011;
				8'b1110010: c <= 9'b1101101;
				8'b1010000: c <= 9'b101001100;
				8'b1111010: c <= 9'b101001;
				8'b1010101: c <= 9'b11110110;
				8'b111011: c <= 9'b100101101;
				8'b1001101: c <= 9'b1;
				8'b111111: c <= 9'b110001011;
				8'b1101110: c <= 9'b101101100;
				8'b1111011: c <= 9'b101110110;
				8'b1001011: c <= 9'b101001100;
				8'b1101111: c <= 9'b1101111;
				8'b1101000: c <= 9'b110100001;
				8'b101100: c <= 9'b11110110;
				8'b100100: c <= 9'b10011001;
				8'b1111000: c <= 9'b101110001;
				8'b1000101: c <= 9'b100111;
				8'b1011001: c <= 9'b101110111;
				8'b110100: c <= 9'b11001100;
				8'b1111001: c <= 9'b10111101;
				8'b1110001: c <= 9'b111000100;
				8'b1001111: c <= 9'b10000;
				8'b1100101: c <= 9'b1000;
				8'b1111110: c <= 9'b101110;
				8'b1111100: c <= 9'b1101100;
				8'b1010110: c <= 9'b100111100;
				8'b110010: c <= 9'b100100101;
				8'b1101101: c <= 9'b10000;
				8'b100011: c <= 9'b111100111;
				8'b1110101: c <= 9'b10111;
				8'b1111101: c <= 9'b101011110;
				8'b101001: c <= 9'b110001100;
				8'b1010010: c <= 9'b101101101;
				8'b1011000: c <= 9'b111100011;
				8'b101110: c <= 9'b110100011;
				8'b1000001: c <= 9'b10010101;
				default: c <= 9'b0;
			endcase
			9'b110111100 : case(di)
				8'b1000011: c <= 9'b100101101;
				8'b101000: c <= 9'b1101001;
				8'b111010: c <= 9'b101110111;
				8'b110110: c <= 9'b100101111;
				8'b1100100: c <= 9'b1011111;
				8'b1000000: c <= 9'b1111;
				8'b1110110: c <= 9'b111011111;
				8'b100101: c <= 9'b11001010;
				8'b101111: c <= 9'b111101000;
				8'b100110: c <= 9'b11100100;
				8'b1100011: c <= 9'b10111101;
				8'b1001000: c <= 9'b100010101;
				8'b111000: c <= 9'b10010000;
				8'b110001: c <= 9'b100100000;
				8'b1010111: c <= 9'b10111100;
				8'b1001110: c <= 9'b100011101;
				8'b1101010: c <= 9'b100110101;
				8'b1001001: c <= 9'b100000010;
				8'b1100000: c <= 9'b111000011;
				8'b110111: c <= 9'b101001100;
				8'b1011101: c <= 9'b111001;
				8'b1011011: c <= 9'b101011101;
				8'b111001: c <= 9'b11111001;
				8'b1001010: c <= 9'b101010100;
				8'b110011: c <= 9'b1000;
				8'b1101100: c <= 9'b11101111;
				8'b1110111: c <= 9'b1111101;
				8'b101011: c <= 9'b11101100;
				8'b1101011: c <= 9'b11111001;
				8'b111100: c <= 9'b100010101;
				8'b1000111: c <= 9'b10111010;
				8'b1011111: c <= 9'b11101;
				8'b1110100: c <= 9'b100010111;
				8'b101101: c <= 9'b100001001;
				8'b1010011: c <= 9'b100101101;
				8'b1100001: c <= 9'b1001001;
				8'b110101: c <= 9'b110000000;
				8'b1000100: c <= 9'b100101111;
				8'b1010001: c <= 9'b110010110;
				8'b1010100: c <= 9'b100000101;
				8'b1100110: c <= 9'b111111011;
				8'b101010: c <= 9'b101111000;
				8'b1011110: c <= 9'b1010111;
				8'b1100111: c <= 9'b1011010;
				8'b1011010: c <= 9'b11111000;
				8'b1000010: c <= 9'b111000000;
				8'b111101: c <= 9'b11010101;
				8'b110000: c <= 9'b111010001;
				8'b111110: c <= 9'b10000001;
				8'b1100010: c <= 9'b111101000;
				8'b1110000: c <= 9'b1101101;
				8'b1101001: c <= 9'b101100000;
				8'b1110011: c <= 9'b100000000;
				8'b1001100: c <= 9'b1000;
				8'b100001: c <= 9'b100010110;
				8'b1000110: c <= 9'b10001011;
				8'b1110010: c <= 9'b1001100;
				8'b1010000: c <= 9'b11111101;
				8'b1111010: c <= 9'b111010;
				8'b1010101: c <= 9'b100110111;
				8'b111011: c <= 9'b101001100;
				8'b1001101: c <= 9'b111001;
				8'b111111: c <= 9'b11000000;
				8'b1101110: c <= 9'b100111001;
				8'b1111011: c <= 9'b1101101;
				8'b1001011: c <= 9'b11100;
				8'b1101111: c <= 9'b110011101;
				8'b1101000: c <= 9'b111111000;
				8'b101100: c <= 9'b111010000;
				8'b100100: c <= 9'b110110101;
				8'b1111000: c <= 9'b100010011;
				8'b1000101: c <= 9'b100100110;
				8'b1011001: c <= 9'b101101001;
				8'b110100: c <= 9'b111110101;
				8'b1111001: c <= 9'b10101110;
				8'b1110001: c <= 9'b10010001;
				8'b1001111: c <= 9'b110001100;
				8'b1100101: c <= 9'b11001110;
				8'b1111110: c <= 9'b100110010;
				8'b1111100: c <= 9'b100001111;
				8'b1010110: c <= 9'b10110001;
				8'b110010: c <= 9'b11100;
				8'b1101101: c <= 9'b10110110;
				8'b100011: c <= 9'b111111001;
				8'b1110101: c <= 9'b101110011;
				8'b1111101: c <= 9'b100101100;
				8'b101001: c <= 9'b10101101;
				8'b1010010: c <= 9'b1111001;
				8'b1011000: c <= 9'b110010011;
				8'b101110: c <= 9'b1001000;
				8'b1000001: c <= 9'b11011010;
				default: c <= 9'b0;
			endcase
			9'b111001010 : case(di)
				8'b1000011: c <= 9'b11011100;
				8'b101000: c <= 9'b11011100;
				8'b111010: c <= 9'b101000110;
				8'b110110: c <= 9'b110010010;
				8'b1100100: c <= 9'b100111;
				8'b1000000: c <= 9'b10000010;
				8'b1110110: c <= 9'b111011100;
				8'b100101: c <= 9'b11010010;
				8'b101111: c <= 9'b111011011;
				8'b100110: c <= 9'b101110;
				8'b1100011: c <= 9'b1110000;
				8'b1001000: c <= 9'b10000110;
				8'b111000: c <= 9'b111111011;
				8'b110001: c <= 9'b1000110;
				8'b1010111: c <= 9'b11110110;
				8'b1001110: c <= 9'b10011100;
				8'b1101010: c <= 9'b101010011;
				8'b1001001: c <= 9'b10000001;
				8'b1100000: c <= 9'b110101101;
				8'b110111: c <= 9'b10100000;
				8'b1011101: c <= 9'b100;
				8'b1011011: c <= 9'b100011001;
				8'b111001: c <= 9'b1111011;
				8'b1001010: c <= 9'b101000010;
				8'b110011: c <= 9'b1000110;
				8'b1101100: c <= 9'b100010;
				8'b1110111: c <= 9'b11010;
				8'b101011: c <= 9'b110010101;
				8'b1101011: c <= 9'b11110100;
				8'b111100: c <= 9'b11111100;
				8'b1000111: c <= 9'b10001111;
				8'b1011111: c <= 9'b100110000;
				8'b1110100: c <= 9'b11001111;
				8'b101101: c <= 9'b11110101;
				8'b1010011: c <= 9'b100000110;
				8'b1100001: c <= 9'b101101;
				8'b110101: c <= 9'b10110110;
				8'b1000100: c <= 9'b111110110;
				8'b1010001: c <= 9'b10010100;
				8'b1010100: c <= 9'b1000111;
				8'b1100110: c <= 9'b101111000;
				8'b101010: c <= 9'b101011;
				8'b1011110: c <= 9'b1000;
				8'b1100111: c <= 9'b1110101;
				8'b1011010: c <= 9'b101010110;
				8'b1000010: c <= 9'b101110101;
				8'b111101: c <= 9'b110110011;
				8'b110000: c <= 9'b101000001;
				8'b111110: c <= 9'b10111100;
				8'b1100010: c <= 9'b110111111;
				8'b1110000: c <= 9'b111001101;
				8'b1101001: c <= 9'b110101100;
				8'b1110011: c <= 9'b1100010;
				8'b1001100: c <= 9'b101100110;
				8'b100001: c <= 9'b111010010;
				8'b1000110: c <= 9'b1111110;
				8'b1110010: c <= 9'b1100;
				8'b1010000: c <= 9'b11000;
				8'b1111010: c <= 9'b1011001;
				8'b1010101: c <= 9'b11111000;
				8'b111011: c <= 9'b110001110;
				8'b1001101: c <= 9'b1001011;
				8'b111111: c <= 9'b110011011;
				8'b1101110: c <= 9'b110100000;
				8'b1111011: c <= 9'b1001000;
				8'b1001011: c <= 9'b110101;
				8'b1101111: c <= 9'b101001001;
				8'b1101000: c <= 9'b101111001;
				8'b101100: c <= 9'b111110000;
				8'b100100: c <= 9'b100000100;
				8'b1111000: c <= 9'b1111100;
				8'b1000101: c <= 9'b11100011;
				8'b1011001: c <= 9'b11101111;
				8'b110100: c <= 9'b1011010;
				8'b1111001: c <= 9'b101100001;
				8'b1110001: c <= 9'b110100;
				8'b1001111: c <= 9'b110001101;
				8'b1100101: c <= 9'b10111010;
				8'b1111110: c <= 9'b110111110;
				8'b1111100: c <= 9'b1111101;
				8'b1010110: c <= 9'b1100011;
				8'b110010: c <= 9'b101110;
				8'b1101101: c <= 9'b1010001;
				8'b100011: c <= 9'b1100111;
				8'b1110101: c <= 9'b1011111;
				8'b1111101: c <= 9'b1000000;
				8'b101001: c <= 9'b10011010;
				8'b1010010: c <= 9'b11100011;
				8'b1011000: c <= 9'b11111100;
				8'b101110: c <= 9'b111101010;
				8'b1000001: c <= 9'b101001000;
				default: c <= 9'b0;
			endcase
			9'b110111001 : case(di)
				8'b1000011: c <= 9'b110011001;
				8'b101000: c <= 9'b100000100;
				8'b111010: c <= 9'b101010011;
				8'b110110: c <= 9'b100000011;
				8'b1100100: c <= 9'b110110000;
				8'b1000000: c <= 9'b101110010;
				8'b1110110: c <= 9'b10101011;
				8'b100101: c <= 9'b1001;
				8'b101111: c <= 9'b110111100;
				8'b100110: c <= 9'b10110101;
				8'b1100011: c <= 9'b111110001;
				8'b1001000: c <= 9'b111101101;
				8'b111000: c <= 9'b1100;
				8'b110001: c <= 9'b110101101;
				8'b1010111: c <= 9'b1010001;
				8'b1001110: c <= 9'b111000000;
				8'b1101010: c <= 9'b111011110;
				8'b1001001: c <= 9'b1110001;
				8'b1100000: c <= 9'b111100001;
				8'b110111: c <= 9'b1101110;
				8'b1011101: c <= 9'b11001101;
				8'b1011011: c <= 9'b100011;
				8'b111001: c <= 9'b100101011;
				8'b1001010: c <= 9'b101110010;
				8'b110011: c <= 9'b11011110;
				8'b1101100: c <= 9'b10001111;
				8'b1110111: c <= 9'b100011010;
				8'b101011: c <= 9'b1001100;
				8'b1101011: c <= 9'b11010101;
				8'b111100: c <= 9'b11100001;
				8'b1000111: c <= 9'b11010111;
				8'b1011111: c <= 9'b111011111;
				8'b1110100: c <= 9'b10010001;
				8'b101101: c <= 9'b11111000;
				8'b1010011: c <= 9'b11010;
				8'b1100001: c <= 9'b111111010;
				8'b110101: c <= 9'b100001111;
				8'b1000100: c <= 9'b111000101;
				8'b1010001: c <= 9'b100110100;
				8'b1010100: c <= 9'b10011011;
				8'b1100110: c <= 9'b1001001;
				8'b101010: c <= 9'b100100011;
				8'b1011110: c <= 9'b11100111;
				8'b1100111: c <= 9'b11011101;
				8'b1011010: c <= 9'b11100111;
				8'b1000010: c <= 9'b110110100;
				8'b111101: c <= 9'b111001111;
				8'b110000: c <= 9'b100110011;
				8'b111110: c <= 9'b100010101;
				8'b1100010: c <= 9'b110010101;
				8'b1110000: c <= 9'b110101011;
				8'b1101001: c <= 9'b110100010;
				8'b1110011: c <= 9'b11100111;
				8'b1001100: c <= 9'b11101011;
				8'b100001: c <= 9'b111000110;
				8'b1000110: c <= 9'b10000111;
				8'b1110010: c <= 9'b111001101;
				8'b1010000: c <= 9'b111010001;
				8'b1111010: c <= 9'b100111101;
				8'b1010101: c <= 9'b11100000;
				8'b111011: c <= 9'b101000101;
				8'b1001101: c <= 9'b11011000;
				8'b111111: c <= 9'b101110100;
				8'b1101110: c <= 9'b11110001;
				8'b1111011: c <= 9'b110100100;
				8'b1001011: c <= 9'b110011011;
				8'b1101111: c <= 9'b101001010;
				8'b1101000: c <= 9'b11111001;
				8'b101100: c <= 9'b10100010;
				8'b100100: c <= 9'b101011110;
				8'b1111000: c <= 9'b100000010;
				8'b1000101: c <= 9'b11110;
				8'b1011001: c <= 9'b101101100;
				8'b110100: c <= 9'b110000;
				8'b1111001: c <= 9'b111000110;
				8'b1110001: c <= 9'b1010001;
				8'b1001111: c <= 9'b10110001;
				8'b1100101: c <= 9'b10001011;
				8'b1111110: c <= 9'b111100101;
				8'b1111100: c <= 9'b100110101;
				8'b1010110: c <= 9'b11111;
				8'b110010: c <= 9'b1111110;
				8'b1101101: c <= 9'b10111101;
				8'b100011: c <= 9'b110110011;
				8'b1110101: c <= 9'b11011100;
				8'b1111101: c <= 9'b10100111;
				8'b101001: c <= 9'b1001010;
				8'b1010010: c <= 9'b10100101;
				8'b1011000: c <= 9'b1011011;
				8'b101110: c <= 9'b100110100;
				8'b1000001: c <= 9'b11010101;
				default: c <= 9'b0;
			endcase
			9'b111101101 : case(di)
				8'b1000011: c <= 9'b101110;
				8'b101000: c <= 9'b101011010;
				8'b111010: c <= 9'b11100101;
				8'b110110: c <= 9'b110101011;
				8'b1100100: c <= 9'b111101010;
				8'b1000000: c <= 9'b101011010;
				8'b1110110: c <= 9'b110100100;
				8'b100101: c <= 9'b10011011;
				8'b101111: c <= 9'b101101001;
				8'b100110: c <= 9'b10011101;
				8'b1100011: c <= 9'b1111111;
				8'b1001000: c <= 9'b10101;
				8'b111000: c <= 9'b100100010;
				8'b110001: c <= 9'b1010110;
				8'b1010111: c <= 9'b101100111;
				8'b1001110: c <= 9'b101100001;
				8'b1101010: c <= 9'b110111100;
				8'b1001001: c <= 9'b110101110;
				8'b1100000: c <= 9'b101110101;
				8'b110111: c <= 9'b110111000;
				8'b1011101: c <= 9'b10101110;
				8'b1011011: c <= 9'b100101100;
				8'b111001: c <= 9'b110111;
				8'b1001010: c <= 9'b111101;
				8'b110011: c <= 9'b1011110;
				8'b1101100: c <= 9'b101010;
				8'b1110111: c <= 9'b10001011;
				8'b101011: c <= 9'b1100000;
				8'b1101011: c <= 9'b100001011;
				8'b111100: c <= 9'b100010110;
				8'b1000111: c <= 9'b100111011;
				8'b1011111: c <= 9'b10110010;
				8'b1110100: c <= 9'b111100100;
				8'b101101: c <= 9'b1001100;
				8'b1010011: c <= 9'b110100100;
				8'b1100001: c <= 9'b111010111;
				8'b110101: c <= 9'b101110010;
				8'b1000100: c <= 9'b101110010;
				8'b1010001: c <= 9'b100111111;
				8'b1010100: c <= 9'b111010100;
				8'b1100110: c <= 9'b110110100;
				8'b101010: c <= 9'b100100001;
				8'b1011110: c <= 9'b10110001;
				8'b1100111: c <= 9'b101110100;
				8'b1011010: c <= 9'b10001111;
				8'b1000010: c <= 9'b110110010;
				8'b111101: c <= 9'b10010;
				8'b110000: c <= 9'b10011011;
				8'b111110: c <= 9'b11010000;
				8'b1100010: c <= 9'b10011000;
				8'b1110000: c <= 9'b100110010;
				8'b1101001: c <= 9'b101010100;
				8'b1110011: c <= 9'b1011;
				8'b1001100: c <= 9'b100011011;
				8'b100001: c <= 9'b111111101;
				8'b1000110: c <= 9'b10111001;
				8'b1110010: c <= 9'b10011100;
				8'b1010000: c <= 9'b111101000;
				8'b1111010: c <= 9'b100110110;
				8'b1010101: c <= 9'b100011011;
				8'b111011: c <= 9'b110111001;
				8'b1001101: c <= 9'b10110110;
				8'b111111: c <= 9'b1010101;
				8'b1101110: c <= 9'b1110000;
				8'b1111011: c <= 9'b110001110;
				8'b1001011: c <= 9'b110001;
				8'b1101111: c <= 9'b101011001;
				8'b1101000: c <= 9'b111110101;
				8'b101100: c <= 9'b11000001;
				8'b100100: c <= 9'b11110111;
				8'b1111000: c <= 9'b110010100;
				8'b1000101: c <= 9'b1011001;
				8'b1011001: c <= 9'b100111001;
				8'b110100: c <= 9'b100100000;
				8'b1111001: c <= 9'b100001010;
				8'b1110001: c <= 9'b10000101;
				8'b1001111: c <= 9'b11000001;
				8'b1100101: c <= 9'b101101000;
				8'b1111110: c <= 9'b101110001;
				8'b1111100: c <= 9'b100001010;
				8'b1010110: c <= 9'b1101100;
				8'b110010: c <= 9'b11111001;
				8'b1101101: c <= 9'b1010001;
				8'b100011: c <= 9'b1001010;
				8'b1110101: c <= 9'b100100000;
				8'b1111101: c <= 9'b100101;
				8'b101001: c <= 9'b110011001;
				8'b1010010: c <= 9'b10010011;
				8'b1011000: c <= 9'b101101010;
				8'b101110: c <= 9'b110001000;
				8'b1000001: c <= 9'b100100010;
				default: c <= 9'b0;
			endcase
			9'b111110110 : case(di)
				8'b1000011: c <= 9'b100010010;
				8'b101000: c <= 9'b11101000;
				8'b111010: c <= 9'b111111101;
				8'b110110: c <= 9'b11011110;
				8'b1100100: c <= 9'b101010000;
				8'b1000000: c <= 9'b10100100;
				8'b1110110: c <= 9'b110111001;
				8'b100101: c <= 9'b11110;
				8'b101111: c <= 9'b111111001;
				8'b100110: c <= 9'b1100100;
				8'b1100011: c <= 9'b11000000;
				8'b1001000: c <= 9'b110101010;
				8'b111000: c <= 9'b110100110;
				8'b110001: c <= 9'b100100101;
				8'b1010111: c <= 9'b101110111;
				8'b1001110: c <= 9'b100101011;
				8'b1101010: c <= 9'b100101110;
				8'b1001001: c <= 9'b1100110;
				8'b1100000: c <= 9'b11001;
				8'b110111: c <= 9'b1100001;
				8'b1011101: c <= 9'b1001001;
				8'b1011011: c <= 9'b111100111;
				8'b111001: c <= 9'b100000111;
				8'b1001010: c <= 9'b11011100;
				8'b110011: c <= 9'b110111111;
				8'b1101100: c <= 9'b11001000;
				8'b1110111: c <= 9'b11110011;
				8'b101011: c <= 9'b111100100;
				8'b1101011: c <= 9'b11011100;
				8'b111100: c <= 9'b101001110;
				8'b1000111: c <= 9'b111010;
				8'b1011111: c <= 9'b110101010;
				8'b1110100: c <= 9'b101111111;
				8'b101101: c <= 9'b100110101;
				8'b1010011: c <= 9'b10111;
				8'b1100001: c <= 9'b1011100;
				8'b110101: c <= 9'b10000101;
				8'b1000100: c <= 9'b100011101;
				8'b1010001: c <= 9'b110000;
				8'b1010100: c <= 9'b110110101;
				8'b1100110: c <= 9'b110100000;
				8'b101010: c <= 9'b11110;
				8'b1011110: c <= 9'b101010000;
				8'b1100111: c <= 9'b110000;
				8'b1011010: c <= 9'b101100000;
				8'b1000010: c <= 9'b100001001;
				8'b111101: c <= 9'b110101101;
				8'b110000: c <= 9'b100000110;
				8'b111110: c <= 9'b101011010;
				8'b1100010: c <= 9'b1110011;
				8'b1110000: c <= 9'b10111000;
				8'b1101001: c <= 9'b10100;
				8'b1110011: c <= 9'b111111000;
				8'b1001100: c <= 9'b100101011;
				8'b100001: c <= 9'b110100;
				8'b1000110: c <= 9'b101110;
				8'b1110010: c <= 9'b110001111;
				8'b1010000: c <= 9'b111001;
				8'b1111010: c <= 9'b11000000;
				8'b1010101: c <= 9'b111001100;
				8'b111011: c <= 9'b110000111;
				8'b1001101: c <= 9'b100111000;
				8'b111111: c <= 9'b101010101;
				8'b1101110: c <= 9'b10011011;
				8'b1111011: c <= 9'b11110000;
				8'b1001011: c <= 9'b111110101;
				8'b1101111: c <= 9'b10110001;
				8'b1101000: c <= 9'b100011010;
				8'b101100: c <= 9'b10010011;
				8'b100100: c <= 9'b110000101;
				8'b1111000: c <= 9'b110111010;
				8'b1000101: c <= 9'b111100011;
				8'b1011001: c <= 9'b111010010;
				8'b110100: c <= 9'b100101111;
				8'b1111001: c <= 9'b11000011;
				8'b1110001: c <= 9'b10010110;
				8'b1001111: c <= 9'b101010;
				8'b1100101: c <= 9'b110100001;
				8'b1111110: c <= 9'b110111011;
				8'b1111100: c <= 9'b101010000;
				8'b1010110: c <= 9'b100110011;
				8'b110010: c <= 9'b101010000;
				8'b1101101: c <= 9'b10000110;
				8'b100011: c <= 9'b1001100;
				8'b1110101: c <= 9'b1001110;
				8'b1111101: c <= 9'b1100010;
				8'b101001: c <= 9'b100000100;
				8'b1010010: c <= 9'b111101001;
				8'b1011000: c <= 9'b100100110;
				8'b101110: c <= 9'b1;
				8'b1000001: c <= 9'b100001001;
				default: c <= 9'b0;
			endcase
			9'b110110000 : case(di)
				8'b1000011: c <= 9'b1110011;
				8'b101000: c <= 9'b1001011;
				8'b111010: c <= 9'b101101110;
				8'b110110: c <= 9'b10100010;
				8'b1100100: c <= 9'b10000111;
				8'b1000000: c <= 9'b10011;
				8'b1110110: c <= 9'b101110011;
				8'b100101: c <= 9'b1010000;
				8'b101111: c <= 9'b10000000;
				8'b100110: c <= 9'b101011101;
				8'b1100011: c <= 9'b100101000;
				8'b1001000: c <= 9'b101100010;
				8'b111000: c <= 9'b101110111;
				8'b110001: c <= 9'b11110;
				8'b1010111: c <= 9'b111000100;
				8'b1001110: c <= 9'b100010010;
				8'b1101010: c <= 9'b101100011;
				8'b1001001: c <= 9'b100011010;
				8'b1100000: c <= 9'b110111001;
				8'b110111: c <= 9'b111010001;
				8'b1011101: c <= 9'b10101001;
				8'b1011011: c <= 9'b1111010;
				8'b111001: c <= 9'b11000000;
				8'b1001010: c <= 9'b101110000;
				8'b110011: c <= 9'b11000100;
				8'b1101100: c <= 9'b110100011;
				8'b1110111: c <= 9'b111111;
				8'b101011: c <= 9'b101001000;
				8'b1101011: c <= 9'b111000100;
				8'b111100: c <= 9'b101111110;
				8'b1000111: c <= 9'b101010110;
				8'b1011111: c <= 9'b10000110;
				8'b1110100: c <= 9'b100100;
				8'b101101: c <= 9'b111101001;
				8'b1010011: c <= 9'b111011110;
				8'b1100001: c <= 9'b11011011;
				8'b110101: c <= 9'b10110100;
				8'b1000100: c <= 9'b1001101;
				8'b1010001: c <= 9'b111100001;
				8'b1010100: c <= 9'b100;
				8'b1100110: c <= 9'b100100001;
				8'b101010: c <= 9'b100100000;
				8'b1011110: c <= 9'b100011100;
				8'b1100111: c <= 9'b11010;
				8'b1011010: c <= 9'b110000;
				8'b1000010: c <= 9'b11100100;
				8'b111101: c <= 9'b100100110;
				8'b110000: c <= 9'b111001011;
				8'b111110: c <= 9'b101001000;
				8'b1100010: c <= 9'b11011;
				8'b1110000: c <= 9'b100101010;
				8'b1101001: c <= 9'b101111010;
				8'b1110011: c <= 9'b110101010;
				8'b1001100: c <= 9'b111000010;
				8'b100001: c <= 9'b11001000;
				8'b1000110: c <= 9'b110010100;
				8'b1110010: c <= 9'b101110010;
				8'b1010000: c <= 9'b10111010;
				8'b1111010: c <= 9'b101111001;
				8'b1010101: c <= 9'b11110011;
				8'b111011: c <= 9'b111111;
				8'b1001101: c <= 9'b10010001;
				8'b111111: c <= 9'b110000011;
				8'b1101110: c <= 9'b100110;
				8'b1111011: c <= 9'b101100000;
				8'b1001011: c <= 9'b111100110;
				8'b1101111: c <= 9'b100101110;
				8'b1101000: c <= 9'b1111110;
				8'b101100: c <= 9'b10111011;
				8'b100100: c <= 9'b101010010;
				8'b1111000: c <= 9'b10101000;
				8'b1000101: c <= 9'b111111001;
				8'b1011001: c <= 9'b101010010;
				8'b110100: c <= 9'b101010000;
				8'b1111001: c <= 9'b110111010;
				8'b1110001: c <= 9'b1011000;
				8'b1001111: c <= 9'b11110000;
				8'b1100101: c <= 9'b11110111;
				8'b1111110: c <= 9'b111001100;
				8'b1111100: c <= 9'b11001100;
				8'b1010110: c <= 9'b111001110;
				8'b110010: c <= 9'b111010010;
				8'b1101101: c <= 9'b1110011;
				8'b100011: c <= 9'b101100001;
				8'b1110101: c <= 9'b10010110;
				8'b1111101: c <= 9'b10101001;
				8'b101001: c <= 9'b100111101;
				8'b1010010: c <= 9'b100111000;
				8'b1011000: c <= 9'b11110000;
				8'b101110: c <= 9'b1100111;
				8'b1000001: c <= 9'b101101101;
				default: c <= 9'b0;
			endcase
			9'b101001 : case(di)
				8'b1000011: c <= 9'b10011101;
				8'b101000: c <= 9'b110111100;
				8'b111010: c <= 9'b1100111;
				8'b110110: c <= 9'b100001100;
				8'b1100100: c <= 9'b1111110;
				8'b1000000: c <= 9'b11011001;
				8'b1110110: c <= 9'b1001101;
				8'b100101: c <= 9'b101010000;
				8'b101111: c <= 9'b1101100;
				8'b100110: c <= 9'b111001110;
				8'b1100011: c <= 9'b101011000;
				8'b1001000: c <= 9'b100000010;
				8'b111000: c <= 9'b1001001;
				8'b110001: c <= 9'b100011;
				8'b1010111: c <= 9'b101010101;
				8'b1001110: c <= 9'b11000011;
				8'b1101010: c <= 9'b11110010;
				8'b1001001: c <= 9'b110000110;
				8'b1100000: c <= 9'b110110000;
				8'b110111: c <= 9'b111010010;
				8'b1011101: c <= 9'b10011111;
				8'b1011011: c <= 9'b1011011;
				8'b111001: c <= 9'b100100110;
				8'b1001010: c <= 9'b1011010;
				8'b110011: c <= 9'b100010100;
				8'b1101100: c <= 9'b110111010;
				8'b1110111: c <= 9'b110001100;
				8'b101011: c <= 9'b110010111;
				8'b1101011: c <= 9'b10101100;
				8'b111100: c <= 9'b101011;
				8'b1000111: c <= 9'b11110001;
				8'b1011111: c <= 9'b11000011;
				8'b1110100: c <= 9'b111001001;
				8'b101101: c <= 9'b11000100;
				8'b1010011: c <= 9'b1100000;
				8'b1100001: c <= 9'b101000101;
				8'b110101: c <= 9'b110111;
				8'b1000100: c <= 9'b1101100;
				8'b1010001: c <= 9'b1000;
				8'b1010100: c <= 9'b111101000;
				8'b1100110: c <= 9'b100010001;
				8'b101010: c <= 9'b1011011;
				8'b1011110: c <= 9'b111101010;
				8'b1100111: c <= 9'b1110000;
				8'b1011010: c <= 9'b10000001;
				8'b1000010: c <= 9'b110111;
				8'b111101: c <= 9'b1101010;
				8'b110000: c <= 9'b110011011;
				8'b111110: c <= 9'b101100110;
				8'b1100010: c <= 9'b10000101;
				8'b1110000: c <= 9'b110011011;
				8'b1101001: c <= 9'b1001110;
				8'b1110011: c <= 9'b100001001;
				8'b1001100: c <= 9'b10001001;
				8'b100001: c <= 9'b111001001;
				8'b1000110: c <= 9'b100010110;
				8'b1110010: c <= 9'b11110011;
				8'b1010000: c <= 9'b1111001;
				8'b1111010: c <= 9'b101100010;
				8'b1010101: c <= 9'b11111101;
				8'b111011: c <= 9'b110001010;
				8'b1001101: c <= 9'b10111111;
				8'b111111: c <= 9'b10011001;
				8'b1101110: c <= 9'b110011010;
				8'b1111011: c <= 9'b100001110;
				8'b1001011: c <= 9'b100110011;
				8'b1101111: c <= 9'b100011100;
				8'b1101000: c <= 9'b101101111;
				8'b101100: c <= 9'b111101100;
				8'b100100: c <= 9'b110110101;
				8'b1111000: c <= 9'b110110;
				8'b1000101: c <= 9'b110000101;
				8'b1011001: c <= 9'b101101110;
				8'b110100: c <= 9'b11110010;
				8'b1111001: c <= 9'b10111101;
				8'b1110001: c <= 9'b100010;
				8'b1001111: c <= 9'b11100001;
				8'b1100101: c <= 9'b11101;
				8'b1111110: c <= 9'b10001100;
				8'b1111100: c <= 9'b1111101;
				8'b1010110: c <= 9'b10010110;
				8'b110010: c <= 9'b111111110;
				8'b1101101: c <= 9'b101000001;
				8'b100011: c <= 9'b10010;
				8'b1110101: c <= 9'b111100001;
				8'b1111101: c <= 9'b110000101;
				8'b101001: c <= 9'b110011101;
				8'b1010010: c <= 9'b110110111;
				8'b1011000: c <= 9'b101100;
				8'b101110: c <= 9'b1000101;
				8'b1000001: c <= 9'b100101110;
				default: c <= 9'b0;
			endcase
			9'b1010001 : case(di)
				8'b1000011: c <= 9'b110001001;
				8'b101000: c <= 9'b111000110;
				8'b111010: c <= 9'b1001101;
				8'b110110: c <= 9'b101101100;
				8'b1100100: c <= 9'b111111000;
				8'b1000000: c <= 9'b11101100;
				8'b1110110: c <= 9'b11001;
				8'b100101: c <= 9'b100011100;
				8'b101111: c <= 9'b1110010;
				8'b100110: c <= 9'b1001110;
				8'b1100011: c <= 9'b1010111;
				8'b1001000: c <= 9'b10010;
				8'b111000: c <= 9'b111001110;
				8'b110001: c <= 9'b11111110;
				8'b1010111: c <= 9'b11100100;
				8'b1001110: c <= 9'b1110101;
				8'b1101010: c <= 9'b101010011;
				8'b1001001: c <= 9'b1111000;
				8'b1100000: c <= 9'b1110101;
				8'b110111: c <= 9'b100110111;
				8'b1011101: c <= 9'b101000011;
				8'b1011011: c <= 9'b111000011;
				8'b111001: c <= 9'b100000101;
				8'b1001010: c <= 9'b111111001;
				8'b110011: c <= 9'b101000;
				8'b1101100: c <= 9'b111100000;
				8'b1110111: c <= 9'b101100101;
				8'b101011: c <= 9'b1010101;
				8'b1101011: c <= 9'b11110000;
				8'b111100: c <= 9'b110001010;
				8'b1000111: c <= 9'b1101101;
				8'b1011111: c <= 9'b110111110;
				8'b1110100: c <= 9'b11011;
				8'b101101: c <= 9'b100010011;
				8'b1010011: c <= 9'b11000011;
				8'b1100001: c <= 9'b101011110;
				8'b110101: c <= 9'b100101111;
				8'b1000100: c <= 9'b1100001;
				8'b1010001: c <= 9'b1011110;
				8'b1010100: c <= 9'b10100100;
				8'b1100110: c <= 9'b110010110;
				8'b101010: c <= 9'b10101011;
				8'b1011110: c <= 9'b11110100;
				8'b1100111: c <= 9'b100100010;
				8'b1011010: c <= 9'b101110100;
				8'b1000010: c <= 9'b10101010;
				8'b111101: c <= 9'b111000010;
				8'b110000: c <= 9'b110001111;
				8'b111110: c <= 9'b111101100;
				8'b1100010: c <= 9'b110101011;
				8'b1110000: c <= 9'b11101011;
				8'b1101001: c <= 9'b110010010;
				8'b1110011: c <= 9'b10000001;
				8'b1001100: c <= 9'b100111000;
				8'b100001: c <= 9'b10000001;
				8'b1000110: c <= 9'b110110101;
				8'b1110010: c <= 9'b101010000;
				8'b1010000: c <= 9'b111111011;
				8'b1111010: c <= 9'b10000111;
				8'b1010101: c <= 9'b110;
				8'b111011: c <= 9'b11110011;
				8'b1001101: c <= 9'b100010111;
				8'b111111: c <= 9'b111001101;
				8'b1101110: c <= 9'b101100110;
				8'b1111011: c <= 9'b110010010;
				8'b1001011: c <= 9'b110111011;
				8'b1101111: c <= 9'b10110011;
				8'b1101000: c <= 9'b110101010;
				8'b101100: c <= 9'b10000001;
				8'b100100: c <= 9'b1001001;
				8'b1111000: c <= 9'b1111111;
				8'b1000101: c <= 9'b10111001;
				8'b1011001: c <= 9'b110001001;
				8'b110100: c <= 9'b100001100;
				8'b1111001: c <= 9'b101110100;
				8'b1110001: c <= 9'b10111011;
				8'b1001111: c <= 9'b100101010;
				8'b1100101: c <= 9'b11000011;
				8'b1111110: c <= 9'b10001011;
				8'b1111100: c <= 9'b10101111;
				8'b1010110: c <= 9'b100000100;
				8'b110010: c <= 9'b101101000;
				8'b1101101: c <= 9'b110000000;
				8'b100011: c <= 9'b111001111;
				8'b1110101: c <= 9'b1100010;
				8'b1111101: c <= 9'b101110011;
				8'b101001: c <= 9'b101101010;
				8'b1010010: c <= 9'b101001111;
				8'b1011000: c <= 9'b111011110;
				8'b101110: c <= 9'b10110010;
				8'b1000001: c <= 9'b111100010;
				default: c <= 9'b0;
			endcase
			9'b111100000 : case(di)
				8'b1000011: c <= 9'b1000011;
				8'b101000: c <= 9'b11101101;
				8'b111010: c <= 9'b1001100;
				8'b110110: c <= 9'b11001111;
				8'b1100100: c <= 9'b1110000;
				8'b1000000: c <= 9'b101111000;
				8'b1110110: c <= 9'b1101001;
				8'b100101: c <= 9'b110001111;
				8'b101111: c <= 9'b10010110;
				8'b100110: c <= 9'b10110100;
				8'b1100011: c <= 9'b11100111;
				8'b1001000: c <= 9'b11000011;
				8'b111000: c <= 9'b101001011;
				8'b110001: c <= 9'b100010010;
				8'b1010111: c <= 9'b11001001;
				8'b1001110: c <= 9'b10000011;
				8'b1101010: c <= 9'b101101101;
				8'b1001001: c <= 9'b110110011;
				8'b1100000: c <= 9'b101011101;
				8'b110111: c <= 9'b10001111;
				8'b1011101: c <= 9'b10110001;
				8'b1011011: c <= 9'b10000001;
				8'b111001: c <= 9'b100111010;
				8'b1001010: c <= 9'b1001110;
				8'b110011: c <= 9'b1011111;
				8'b1101100: c <= 9'b10101101;
				8'b1110111: c <= 9'b11110110;
				8'b101011: c <= 9'b111100;
				8'b1101011: c <= 9'b101001000;
				8'b111100: c <= 9'b111101101;
				8'b1000111: c <= 9'b101010100;
				8'b1011111: c <= 9'b100000001;
				8'b1110100: c <= 9'b11011000;
				8'b101101: c <= 9'b111010;
				8'b1010011: c <= 9'b101111000;
				8'b1100001: c <= 9'b1110010;
				8'b110101: c <= 9'b1000011;
				8'b1000100: c <= 9'b1010010;
				8'b1010001: c <= 9'b111111101;
				8'b1010100: c <= 9'b110100010;
				8'b1100110: c <= 9'b100011101;
				8'b101010: c <= 9'b11100001;
				8'b1011110: c <= 9'b1111100;
				8'b1100111: c <= 9'b10111001;
				8'b1011010: c <= 9'b110010110;
				8'b1000010: c <= 9'b10010;
				8'b111101: c <= 9'b1111000;
				8'b110000: c <= 9'b1011010;
				8'b111110: c <= 9'b111100000;
				8'b1100010: c <= 9'b111101110;
				8'b1110000: c <= 9'b1000111;
				8'b1101001: c <= 9'b10011010;
				8'b1110011: c <= 9'b100010110;
				8'b1001100: c <= 9'b1101010;
				8'b100001: c <= 9'b110010001;
				8'b1000110: c <= 9'b11010;
				8'b1110010: c <= 9'b101111000;
				8'b1010000: c <= 9'b110000011;
				8'b1111010: c <= 9'b1000010;
				8'b1010101: c <= 9'b1001111;
				8'b111011: c <= 9'b11110100;
				8'b1001101: c <= 9'b1001;
				8'b111111: c <= 9'b111001001;
				8'b1101110: c <= 9'b10111111;
				8'b1111011: c <= 9'b11010000;
				8'b1001011: c <= 9'b100101110;
				8'b1101111: c <= 9'b1100001;
				8'b1101000: c <= 9'b100101000;
				8'b101100: c <= 9'b111001011;
				8'b100100: c <= 9'b110111110;
				8'b1111000: c <= 9'b100100001;
				8'b1000101: c <= 9'b110100111;
				8'b1011001: c <= 9'b1111111;
				8'b110100: c <= 9'b110001011;
				8'b1111001: c <= 9'b101111010;
				8'b1110001: c <= 9'b11100111;
				8'b1001111: c <= 9'b111110110;
				8'b1100101: c <= 9'b100001;
				8'b1111110: c <= 9'b1101000;
				8'b1111100: c <= 9'b111110000;
				8'b1010110: c <= 9'b101100011;
				8'b110010: c <= 9'b111000011;
				8'b1101101: c <= 9'b100101;
				8'b100011: c <= 9'b101010110;
				8'b1110101: c <= 9'b10010111;
				8'b1111101: c <= 9'b10101111;
				8'b101001: c <= 9'b100010;
				8'b1010010: c <= 9'b111001011;
				8'b1011000: c <= 9'b111101101;
				8'b101110: c <= 9'b101110001;
				8'b1000001: c <= 9'b100110101;
				default: c <= 9'b0;
			endcase
			9'b110010111 : case(di)
				8'b1000011: c <= 9'b101001010;
				8'b101000: c <= 9'b110110010;
				8'b111010: c <= 9'b100010101;
				8'b110110: c <= 9'b101001000;
				8'b1100100: c <= 9'b10000;
				8'b1000000: c <= 9'b101011;
				8'b1110110: c <= 9'b1001;
				8'b100101: c <= 9'b100110010;
				8'b101111: c <= 9'b10101010;
				8'b100110: c <= 9'b10000001;
				8'b1100011: c <= 9'b1100000;
				8'b1001000: c <= 9'b101000111;
				8'b111000: c <= 9'b101101111;
				8'b110001: c <= 9'b1110111;
				8'b1010111: c <= 9'b101010000;
				8'b1001110: c <= 9'b110011111;
				8'b1101010: c <= 9'b11110011;
				8'b1001001: c <= 9'b10001000;
				8'b1100000: c <= 9'b11011101;
				8'b110111: c <= 9'b11011110;
				8'b1011101: c <= 9'b11110111;
				8'b1011011: c <= 9'b110011110;
				8'b111001: c <= 9'b111000011;
				8'b1001010: c <= 9'b10010100;
				8'b110011: c <= 9'b100010000;
				8'b1101100: c <= 9'b111011;
				8'b1110111: c <= 9'b1100001;
				8'b101011: c <= 9'b11001;
				8'b1101011: c <= 9'b1011;
				8'b111100: c <= 9'b10101000;
				8'b1000111: c <= 9'b10010111;
				8'b1011111: c <= 9'b11111001;
				8'b1110100: c <= 9'b10011011;
				8'b101101: c <= 9'b101011110;
				8'b1010011: c <= 9'b10010100;
				8'b1100001: c <= 9'b100111111;
				8'b110101: c <= 9'b110010;
				8'b1000100: c <= 9'b100011111;
				8'b1010001: c <= 9'b11110100;
				8'b1010100: c <= 9'b10110110;
				8'b1100110: c <= 9'b1111;
				8'b101010: c <= 9'b10101010;
				8'b1011110: c <= 9'b10011010;
				8'b1100111: c <= 9'b11011101;
				8'b1011010: c <= 9'b1111010;
				8'b1000010: c <= 9'b111001011;
				8'b111101: c <= 9'b10010001;
				8'b110000: c <= 9'b11101011;
				8'b111110: c <= 9'b111101100;
				8'b1100010: c <= 9'b1011111;
				8'b1110000: c <= 9'b1100101;
				8'b1101001: c <= 9'b110000;
				8'b1110011: c <= 9'b11011110;
				8'b1001100: c <= 9'b101010000;
				8'b100001: c <= 9'b10011010;
				8'b1000110: c <= 9'b10101010;
				8'b1110010: c <= 9'b11101111;
				8'b1010000: c <= 9'b110111011;
				8'b1111010: c <= 9'b101110001;
				8'b1010101: c <= 9'b10000111;
				8'b111011: c <= 9'b100110100;
				8'b1001101: c <= 9'b111001010;
				8'b111111: c <= 9'b111101111;
				8'b1101110: c <= 9'b11110111;
				8'b1111011: c <= 9'b110100001;
				8'b1001011: c <= 9'b10000010;
				8'b1101111: c <= 9'b111001111;
				8'b1101000: c <= 9'b101100001;
				8'b101100: c <= 9'b1011111;
				8'b100100: c <= 9'b100111011;
				8'b1111000: c <= 9'b11011;
				8'b1000101: c <= 9'b10001000;
				8'b1011001: c <= 9'b11100001;
				8'b110100: c <= 9'b11000010;
				8'b1111001: c <= 9'b1000101;
				8'b1110001: c <= 9'b110000010;
				8'b1001111: c <= 9'b111011110;
				8'b1100101: c <= 9'b11010001;
				8'b1111110: c <= 9'b11001001;
				8'b1111100: c <= 9'b101110011;
				8'b1010110: c <= 9'b110011110;
				8'b110010: c <= 9'b1011011;
				8'b1101101: c <= 9'b110101101;
				8'b100011: c <= 9'b100100101;
				8'b1110101: c <= 9'b100011;
				8'b1111101: c <= 9'b110100101;
				8'b101001: c <= 9'b11000010;
				8'b1010010: c <= 9'b101110010;
				8'b1011000: c <= 9'b10010100;
				8'b101110: c <= 9'b111001110;
				8'b1000001: c <= 9'b11101000;
				default: c <= 9'b0;
			endcase
			9'b10101100 : case(di)
				8'b1000011: c <= 9'b111000011;
				8'b101000: c <= 9'b11001100;
				8'b111010: c <= 9'b111110110;
				8'b110110: c <= 9'b101100010;
				8'b1100100: c <= 9'b1111110;
				8'b1000000: c <= 9'b1111110;
				8'b1110110: c <= 9'b11110;
				8'b100101: c <= 9'b110100101;
				8'b101111: c <= 9'b111110001;
				8'b100110: c <= 9'b100;
				8'b1100011: c <= 9'b111111110;
				8'b1001000: c <= 9'b1000110;
				8'b111000: c <= 9'b101101011;
				8'b110001: c <= 9'b1000111;
				8'b1010111: c <= 9'b10000001;
				8'b1001110: c <= 9'b1110010;
				8'b1101010: c <= 9'b11011110;
				8'b1001001: c <= 9'b100110;
				8'b1100000: c <= 9'b110111100;
				8'b110111: c <= 9'b100011011;
				8'b1011101: c <= 9'b110110;
				8'b1011011: c <= 9'b111010100;
				8'b111001: c <= 9'b10011101;
				8'b1001010: c <= 9'b100000100;
				8'b110011: c <= 9'b11011101;
				8'b1101100: c <= 9'b11001111;
				8'b1110111: c <= 9'b110100001;
				8'b101011: c <= 9'b10100000;
				8'b1101011: c <= 9'b11101;
				8'b111100: c <= 9'b1011100;
				8'b1000111: c <= 9'b11101101;
				8'b1011111: c <= 9'b11100001;
				8'b1110100: c <= 9'b100101010;
				8'b101101: c <= 9'b101110010;
				8'b1010011: c <= 9'b111001;
				8'b1100001: c <= 9'b111011001;
				8'b110101: c <= 9'b101111010;
				8'b1000100: c <= 9'b111010000;
				8'b1010001: c <= 9'b110000010;
				8'b1010100: c <= 9'b101101011;
				8'b1100110: c <= 9'b101110110;
				8'b101010: c <= 9'b1100001;
				8'b1011110: c <= 9'b1111100;
				8'b1100111: c <= 9'b111000011;
				8'b1011010: c <= 9'b1001;
				8'b1000010: c <= 9'b10101111;
				8'b111101: c <= 9'b111000100;
				8'b110000: c <= 9'b1101;
				8'b111110: c <= 9'b111111011;
				8'b1100010: c <= 9'b10011100;
				8'b1110000: c <= 9'b111010000;
				8'b1101001: c <= 9'b111;
				8'b1110011: c <= 9'b10101111;
				8'b1001100: c <= 9'b111000010;
				8'b100001: c <= 9'b11000000;
				8'b1000110: c <= 9'b11101000;
				8'b1110010: c <= 9'b10010000;
				8'b1010000: c <= 9'b100101001;
				8'b1111010: c <= 9'b10010;
				8'b1010101: c <= 9'b11011;
				8'b111011: c <= 9'b1101101;
				8'b1001101: c <= 9'b111000010;
				8'b111111: c <= 9'b101110001;
				8'b1101110: c <= 9'b110111;
				8'b1111011: c <= 9'b11000010;
				8'b1001011: c <= 9'b110110011;
				8'b1101111: c <= 9'b100111;
				8'b1101000: c <= 9'b100010100;
				8'b101100: c <= 9'b11011101;
				8'b100100: c <= 9'b1100111;
				8'b1111000: c <= 9'b110101011;
				8'b1000101: c <= 9'b111001010;
				8'b1011001: c <= 9'b1100110;
				8'b110100: c <= 9'b10101;
				8'b1111001: c <= 9'b11011100;
				8'b1110001: c <= 9'b110110101;
				8'b1001111: c <= 9'b101110100;
				8'b1100101: c <= 9'b101011011;
				8'b1111110: c <= 9'b10001001;
				8'b1111100: c <= 9'b1110101;
				8'b1010110: c <= 9'b11100001;
				8'b110010: c <= 9'b110010010;
				8'b1101101: c <= 9'b11001010;
				8'b100011: c <= 9'b11100111;
				8'b1110101: c <= 9'b100101111;
				8'b1111101: c <= 9'b111001100;
				8'b101001: c <= 9'b101001110;
				8'b1010010: c <= 9'b11100011;
				8'b1011000: c <= 9'b101101111;
				8'b101110: c <= 9'b11001110;
				8'b1000001: c <= 9'b100111;
				default: c <= 9'b0;
			endcase
			9'b100000001 : case(di)
				8'b1000011: c <= 9'b11011011;
				8'b101000: c <= 9'b10001101;
				8'b111010: c <= 9'b111001110;
				8'b110110: c <= 9'b101001100;
				8'b1100100: c <= 9'b11110110;
				8'b1000000: c <= 9'b100010011;
				8'b1110110: c <= 9'b100001101;
				8'b100101: c <= 9'b110011;
				8'b101111: c <= 9'b1010010;
				8'b100110: c <= 9'b111100110;
				8'b1100011: c <= 9'b110111;
				8'b1001000: c <= 9'b110011100;
				8'b111000: c <= 9'b100110011;
				8'b110001: c <= 9'b1111110;
				8'b1010111: c <= 9'b110000110;
				8'b1001110: c <= 9'b10100100;
				8'b1101010: c <= 9'b110000111;
				8'b1001001: c <= 9'b101101010;
				8'b1100000: c <= 9'b1110101;
				8'b110111: c <= 9'b11111000;
				8'b1011101: c <= 9'b1000110;
				8'b1011011: c <= 9'b111100100;
				8'b111001: c <= 9'b101111111;
				8'b1001010: c <= 9'b101100011;
				8'b110011: c <= 9'b10110011;
				8'b1101100: c <= 9'b111100011;
				8'b1110111: c <= 9'b101010001;
				8'b101011: c <= 9'b1001;
				8'b1101011: c <= 9'b10010;
				8'b111100: c <= 9'b100;
				8'b1000111: c <= 9'b110001010;
				8'b1011111: c <= 9'b1111;
				8'b1110100: c <= 9'b1;
				8'b101101: c <= 9'b10;
				8'b1010011: c <= 9'b111001010;
				8'b1100001: c <= 9'b11110110;
				8'b110101: c <= 9'b110110101;
				8'b1000100: c <= 9'b111100011;
				8'b1010001: c <= 9'b110011001;
				8'b1010100: c <= 9'b10001111;
				8'b1100110: c <= 9'b101110110;
				8'b101010: c <= 9'b101000011;
				8'b1011110: c <= 9'b110000000;
				8'b1100111: c <= 9'b101101101;
				8'b1011010: c <= 9'b10011100;
				8'b1000010: c <= 9'b101100000;
				8'b111101: c <= 9'b101110;
				8'b110000: c <= 9'b11111010;
				8'b111110: c <= 9'b10111111;
				8'b1100010: c <= 9'b111011110;
				8'b1110000: c <= 9'b101100011;
				8'b1101001: c <= 9'b1101110;
				8'b1110011: c <= 9'b11010100;
				8'b1001100: c <= 9'b110000;
				8'b100001: c <= 9'b11111110;
				8'b1000110: c <= 9'b110001;
				8'b1110010: c <= 9'b111101001;
				8'b1010000: c <= 9'b100101000;
				8'b1111010: c <= 9'b100110101;
				8'b1010101: c <= 9'b11000111;
				8'b111011: c <= 9'b110101110;
				8'b1001101: c <= 9'b1110111;
				8'b111111: c <= 9'b110011111;
				8'b1101110: c <= 9'b111101010;
				8'b1111011: c <= 9'b10101101;
				8'b1001011: c <= 9'b1100;
				8'b1101111: c <= 9'b11000110;
				8'b1101000: c <= 9'b111;
				8'b101100: c <= 9'b1000011;
				8'b100100: c <= 9'b110111010;
				8'b1111000: c <= 9'b10010101;
				8'b1000101: c <= 9'b110010001;
				8'b1011001: c <= 9'b1011001;
				8'b110100: c <= 9'b110100100;
				8'b1111001: c <= 9'b1101000;
				8'b1110001: c <= 9'b11100000;
				8'b1001111: c <= 9'b11011001;
				8'b1100101: c <= 9'b101101;
				8'b1111110: c <= 9'b111110101;
				8'b1111100: c <= 9'b111000101;
				8'b1010110: c <= 9'b110101111;
				8'b110010: c <= 9'b101011;
				8'b1101101: c <= 9'b110100011;
				8'b100011: c <= 9'b10111000;
				8'b1110101: c <= 9'b100111100;
				8'b1111101: c <= 9'b1000;
				8'b101001: c <= 9'b110100111;
				8'b1010010: c <= 9'b10010111;
				8'b1011000: c <= 9'b10011001;
				8'b101110: c <= 9'b101110;
				8'b1000001: c <= 9'b1111001;
				default: c <= 9'b0;
			endcase
			9'b110101010 : case(di)
				8'b1000011: c <= 9'b111000111;
				8'b101000: c <= 9'b101100100;
				8'b111010: c <= 9'b101;
				8'b110110: c <= 9'b111011010;
				8'b1100100: c <= 9'b10111001;
				8'b1000000: c <= 9'b101101001;
				8'b1110110: c <= 9'b111101100;
				8'b100101: c <= 9'b101011010;
				8'b101111: c <= 9'b110010001;
				8'b100110: c <= 9'b101100011;
				8'b1100011: c <= 9'b1111010;
				8'b1001000: c <= 9'b11;
				8'b111000: c <= 9'b11000;
				8'b110001: c <= 9'b110101011;
				8'b1010111: c <= 9'b11011011;
				8'b1001110: c <= 9'b100110;
				8'b1101010: c <= 9'b100010011;
				8'b1001001: c <= 9'b1;
				8'b1100000: c <= 9'b11110111;
				8'b110111: c <= 9'b1000000;
				8'b1011101: c <= 9'b1101010;
				8'b1011011: c <= 9'b10000101;
				8'b111001: c <= 9'b101010100;
				8'b1001010: c <= 9'b11100000;
				8'b110011: c <= 9'b100111101;
				8'b1101100: c <= 9'b111010010;
				8'b1110111: c <= 9'b101110;
				8'b101011: c <= 9'b1001101;
				8'b1101011: c <= 9'b1111111;
				8'b111100: c <= 9'b100100001;
				8'b1000111: c <= 9'b111111;
				8'b1011111: c <= 9'b100101111;
				8'b1110100: c <= 9'b10101011;
				8'b101101: c <= 9'b111000100;
				8'b1010011: c <= 9'b111000010;
				8'b1100001: c <= 9'b1101000;
				8'b110101: c <= 9'b101011101;
				8'b1000100: c <= 9'b1101111;
				8'b1010001: c <= 9'b101010100;
				8'b1010100: c <= 9'b100010110;
				8'b1100110: c <= 9'b110111;
				8'b101010: c <= 9'b1011011;
				8'b1011110: c <= 9'b1011110;
				8'b1100111: c <= 9'b1011001;
				8'b1011010: c <= 9'b101;
				8'b1000010: c <= 9'b100010;
				8'b111101: c <= 9'b111001111;
				8'b110000: c <= 9'b100101011;
				8'b111110: c <= 9'b110101001;
				8'b1100010: c <= 9'b100110100;
				8'b1110000: c <= 9'b111001001;
				8'b1101001: c <= 9'b110111010;
				8'b1110011: c <= 9'b111010000;
				8'b1001100: c <= 9'b1010001;
				8'b100001: c <= 9'b100011101;
				8'b1000110: c <= 9'b10111110;
				8'b1110010: c <= 9'b1001110;
				8'b1010000: c <= 9'b100001;
				8'b1111010: c <= 9'b10011010;
				8'b1010101: c <= 9'b10111010;
				8'b111011: c <= 9'b11111100;
				8'b1001101: c <= 9'b10110111;
				8'b111111: c <= 9'b101111000;
				8'b1101110: c <= 9'b10001011;
				8'b1111011: c <= 9'b100110100;
				8'b1001011: c <= 9'b11001110;
				8'b1101111: c <= 9'b10;
				8'b1101000: c <= 9'b111111001;
				8'b101100: c <= 9'b100101011;
				8'b100100: c <= 9'b1001110;
				8'b1111000: c <= 9'b10000001;
				8'b1000101: c <= 9'b110000;
				8'b1011001: c <= 9'b1000001;
				8'b110100: c <= 9'b1011000;
				8'b1111001: c <= 9'b10100;
				8'b1110001: c <= 9'b100000000;
				8'b1001111: c <= 9'b110010001;
				8'b1100101: c <= 9'b111000;
				8'b1111110: c <= 9'b100100000;
				8'b1111100: c <= 9'b111;
				8'b1010110: c <= 9'b1110010;
				8'b110010: c <= 9'b110101111;
				8'b1101101: c <= 9'b101101110;
				8'b100011: c <= 9'b100110010;
				8'b1110101: c <= 9'b1100001;
				8'b1111101: c <= 9'b111010001;
				8'b101001: c <= 9'b11001010;
				8'b1010010: c <= 9'b111010;
				8'b1011000: c <= 9'b111100001;
				8'b101110: c <= 9'b11100110;
				8'b1000001: c <= 9'b111100011;
				default: c <= 9'b0;
			endcase
			9'b11001000 : case(di)
				8'b1000011: c <= 9'b111000101;
				8'b101000: c <= 9'b10010101;
				8'b111010: c <= 9'b11110010;
				8'b110110: c <= 9'b100001110;
				8'b1100100: c <= 9'b1001001;
				8'b1000000: c <= 9'b111000000;
				8'b1110110: c <= 9'b111011001;
				8'b100101: c <= 9'b111110101;
				8'b101111: c <= 9'b110111011;
				8'b100110: c <= 9'b111010110;
				8'b1100011: c <= 9'b10100;
				8'b1001000: c <= 9'b1001001;
				8'b111000: c <= 9'b1001000;
				8'b110001: c <= 9'b11010111;
				8'b1010111: c <= 9'b1000001;
				8'b1001110: c <= 9'b110011101;
				8'b1101010: c <= 9'b111101000;
				8'b1001001: c <= 9'b101000011;
				8'b1100000: c <= 9'b111011100;
				8'b110111: c <= 9'b11110101;
				8'b1011101: c <= 9'b100110011;
				8'b1011011: c <= 9'b111111010;
				8'b111001: c <= 9'b10101100;
				8'b1001010: c <= 9'b10101100;
				8'b110011: c <= 9'b11111000;
				8'b1101100: c <= 9'b100100001;
				8'b1110111: c <= 9'b100100111;
				8'b101011: c <= 9'b111000011;
				8'b1101011: c <= 9'b11000000;
				8'b111100: c <= 9'b11000010;
				8'b1000111: c <= 9'b111111101;
				8'b1011111: c <= 9'b100;
				8'b1110100: c <= 9'b100110101;
				8'b101101: c <= 9'b11001101;
				8'b1010011: c <= 9'b1101;
				8'b1100001: c <= 9'b11110110;
				8'b110101: c <= 9'b101010;
				8'b1000100: c <= 9'b11100010;
				8'b1010001: c <= 9'b110011100;
				8'b1010100: c <= 9'b110010101;
				8'b1100110: c <= 9'b11110000;
				8'b101010: c <= 9'b101010111;
				8'b1011110: c <= 9'b101001110;
				8'b1100111: c <= 9'b100101111;
				8'b1011010: c <= 9'b101110010;
				8'b1000010: c <= 9'b10100011;
				8'b111101: c <= 9'b1000011;
				8'b110000: c <= 9'b1000110;
				8'b111110: c <= 9'b110111110;
				8'b1100010: c <= 9'b101101011;
				8'b1110000: c <= 9'b1000;
				8'b1101001: c <= 9'b1101;
				8'b1110011: c <= 9'b100110110;
				8'b1001100: c <= 9'b111100;
				8'b100001: c <= 9'b110110111;
				8'b1000110: c <= 9'b10101001;
				8'b1110010: c <= 9'b111100100;
				8'b1010000: c <= 9'b100010110;
				8'b1111010: c <= 9'b101101011;
				8'b1010101: c <= 9'b10111101;
				8'b111011: c <= 9'b10101110;
				8'b1001101: c <= 9'b1001;
				8'b111111: c <= 9'b110010111;
				8'b1101110: c <= 9'b1101110;
				8'b1111011: c <= 9'b101111111;
				8'b1001011: c <= 9'b11000100;
				8'b1101111: c <= 9'b100001111;
				8'b1101000: c <= 9'b101111000;
				8'b101100: c <= 9'b11011011;
				8'b100100: c <= 9'b100011;
				8'b1111000: c <= 9'b111101001;
				8'b1000101: c <= 9'b10100000;
				8'b1011001: c <= 9'b111100100;
				8'b110100: c <= 9'b101010000;
				8'b1111001: c <= 9'b101100111;
				8'b1110001: c <= 9'b111101010;
				8'b1001111: c <= 9'b111100001;
				8'b1100101: c <= 9'b100100110;
				8'b1111110: c <= 9'b1110001;
				8'b1111100: c <= 9'b10011010;
				8'b1010110: c <= 9'b111101000;
				8'b110010: c <= 9'b10100011;
				8'b1101101: c <= 9'b1100100;
				8'b100011: c <= 9'b101110101;
				8'b1110101: c <= 9'b110001001;
				8'b1111101: c <= 9'b101001011;
				8'b101001: c <= 9'b110001;
				8'b1010010: c <= 9'b11011101;
				8'b1011000: c <= 9'b1101101;
				8'b101110: c <= 9'b11111;
				8'b1000001: c <= 9'b111000011;
				default: c <= 9'b0;
			endcase
			9'b101100111 : case(di)
				8'b1000011: c <= 9'b11100011;
				8'b101000: c <= 9'b1010110;
				8'b111010: c <= 9'b1101100;
				8'b110110: c <= 9'b110101001;
				8'b1100100: c <= 9'b100110;
				8'b1000000: c <= 9'b101010000;
				8'b1110110: c <= 9'b101100110;
				8'b100101: c <= 9'b1000001;
				8'b101111: c <= 9'b101001010;
				8'b100110: c <= 9'b100110110;
				8'b1100011: c <= 9'b111000100;
				8'b1001000: c <= 9'b100010000;
				8'b111000: c <= 9'b100111111;
				8'b110001: c <= 9'b11001001;
				8'b1010111: c <= 9'b111010000;
				8'b1001110: c <= 9'b1111001;
				8'b1101010: c <= 9'b11011011;
				8'b1001001: c <= 9'b11011000;
				8'b1100000: c <= 9'b110001;
				8'b110111: c <= 9'b1111011;
				8'b1011101: c <= 9'b101010000;
				8'b1011011: c <= 9'b11110011;
				8'b111001: c <= 9'b111111110;
				8'b1001010: c <= 9'b101001000;
				8'b110011: c <= 9'b100001;
				8'b1101100: c <= 9'b100100010;
				8'b1110111: c <= 9'b110111010;
				8'b101011: c <= 9'b11011101;
				8'b1101011: c <= 9'b111010110;
				8'b111100: c <= 9'b110110100;
				8'b1000111: c <= 9'b110;
				8'b1011111: c <= 9'b101001001;
				8'b1110100: c <= 9'b10001010;
				8'b101101: c <= 9'b110010110;
				8'b1010011: c <= 9'b1100011;
				8'b1100001: c <= 9'b100100111;
				8'b110101: c <= 9'b111011110;
				8'b1000100: c <= 9'b11110001;
				8'b1010001: c <= 9'b110010110;
				8'b1010100: c <= 9'b11001111;
				8'b1100110: c <= 9'b10011111;
				8'b101010: c <= 9'b100011001;
				8'b1011110: c <= 9'b111000111;
				8'b1100111: c <= 9'b100000000;
				8'b1011010: c <= 9'b101011111;
				8'b1000010: c <= 9'b100011;
				8'b111101: c <= 9'b101010000;
				8'b110000: c <= 9'b100100110;
				8'b111110: c <= 9'b11101101;
				8'b1100010: c <= 9'b11111001;
				8'b1110000: c <= 9'b101110;
				8'b1101001: c <= 9'b10110;
				8'b1110011: c <= 9'b1001001;
				8'b1001100: c <= 9'b10010111;
				8'b100001: c <= 9'b10100100;
				8'b1000110: c <= 9'b11101100;
				8'b1110010: c <= 9'b11110;
				8'b1010000: c <= 9'b111101101;
				8'b1111010: c <= 9'b100110010;
				8'b1010101: c <= 9'b1011011;
				8'b111011: c <= 9'b100110110;
				8'b1001101: c <= 9'b110100011;
				8'b111111: c <= 9'b101011010;
				8'b1101110: c <= 9'b111110011;
				8'b1111011: c <= 9'b1011110;
				8'b1001011: c <= 9'b10011010;
				8'b1101111: c <= 9'b11111101;
				8'b1101000: c <= 9'b110101011;
				8'b101100: c <= 9'b111111111;
				8'b100100: c <= 9'b101011111;
				8'b1111000: c <= 9'b10010;
				8'b1000101: c <= 9'b110011100;
				8'b1011001: c <= 9'b10110001;
				8'b110100: c <= 9'b111100000;
				8'b1111001: c <= 9'b110101100;
				8'b1110001: c <= 9'b110011010;
				8'b1001111: c <= 9'b110101001;
				8'b1100101: c <= 9'b100101101;
				8'b1111110: c <= 9'b1001101;
				8'b1111100: c <= 9'b110111000;
				8'b1010110: c <= 9'b100011000;
				8'b110010: c <= 9'b101101101;
				8'b1101101: c <= 9'b10001111;
				8'b100011: c <= 9'b11100000;
				8'b1110101: c <= 9'b11000011;
				8'b1111101: c <= 9'b1001101;
				8'b101001: c <= 9'b100101;
				8'b1010010: c <= 9'b101010110;
				8'b1011000: c <= 9'b111101100;
				8'b101110: c <= 9'b11110011;
				8'b1000001: c <= 9'b10001011;
				default: c <= 9'b0;
			endcase
			9'b10111101 : case(di)
				8'b1000011: c <= 9'b11010010;
				8'b101000: c <= 9'b110101001;
				8'b111010: c <= 9'b111110101;
				8'b110110: c <= 9'b110011111;
				8'b1100100: c <= 9'b100100101;
				8'b1000000: c <= 9'b110;
				8'b1110110: c <= 9'b11000000;
				8'b100101: c <= 9'b101101101;
				8'b101111: c <= 9'b100111000;
				8'b100110: c <= 9'b1011010;
				8'b1100011: c <= 9'b1100101;
				8'b1001000: c <= 9'b100001100;
				8'b111000: c <= 9'b100101010;
				8'b110001: c <= 9'b1111100;
				8'b1010111: c <= 9'b101111110;
				8'b1001110: c <= 9'b100111000;
				8'b1101010: c <= 9'b10001111;
				8'b1001001: c <= 9'b100001001;
				8'b1100000: c <= 9'b1101;
				8'b110111: c <= 9'b110111110;
				8'b1011101: c <= 9'b110101010;
				8'b1011011: c <= 9'b10011100;
				8'b111001: c <= 9'b1010000;
				8'b1001010: c <= 9'b110101010;
				8'b110011: c <= 9'b10100;
				8'b1101100: c <= 9'b1101101;
				8'b1110111: c <= 9'b10101011;
				8'b101011: c <= 9'b101100111;
				8'b1101011: c <= 9'b110111111;
				8'b111100: c <= 9'b101000111;
				8'b1000111: c <= 9'b101011010;
				8'b1011111: c <= 9'b111000010;
				8'b1110100: c <= 9'b100011001;
				8'b101101: c <= 9'b110111111;
				8'b1010011: c <= 9'b1000111;
				8'b1100001: c <= 9'b10110010;
				8'b110101: c <= 9'b100011;
				8'b1000100: c <= 9'b11100110;
				8'b1010001: c <= 9'b1110111;
				8'b1010100: c <= 9'b100111000;
				8'b1100110: c <= 9'b101111010;
				8'b101010: c <= 9'b101000111;
				8'b1011110: c <= 9'b110011100;
				8'b1100111: c <= 9'b111001110;
				8'b1011010: c <= 9'b100100011;
				8'b1000010: c <= 9'b101111001;
				8'b111101: c <= 9'b101011000;
				8'b110000: c <= 9'b1100010;
				8'b111110: c <= 9'b10000110;
				8'b1100010: c <= 9'b10111101;
				8'b1110000: c <= 9'b111001011;
				8'b1101001: c <= 9'b100111000;
				8'b1110011: c <= 9'b110000;
				8'b1001100: c <= 9'b10010;
				8'b100001: c <= 9'b111000100;
				8'b1000110: c <= 9'b11000000;
				8'b1110010: c <= 9'b100110010;
				8'b1010000: c <= 9'b1111011;
				8'b1111010: c <= 9'b100010111;
				8'b1010101: c <= 9'b11001001;
				8'b111011: c <= 9'b1010001;
				8'b1001101: c <= 9'b101100110;
				8'b111111: c <= 9'b100001011;
				8'b1101110: c <= 9'b110110010;
				8'b1111011: c <= 9'b1000101;
				8'b1001011: c <= 9'b10010111;
				8'b1101111: c <= 9'b1001100;
				8'b1101000: c <= 9'b100101011;
				8'b101100: c <= 9'b11001001;
				8'b100100: c <= 9'b101110101;
				8'b1111000: c <= 9'b100001;
				8'b1000101: c <= 9'b110100001;
				8'b1011001: c <= 9'b10001101;
				8'b110100: c <= 9'b111100011;
				8'b1111001: c <= 9'b111010111;
				8'b1110001: c <= 9'b1001110;
				8'b1001111: c <= 9'b111111011;
				8'b1100101: c <= 9'b10001000;
				8'b1111110: c <= 9'b100011100;
				8'b1111100: c <= 9'b100111111;
				8'b1010110: c <= 9'b111100100;
				8'b110010: c <= 9'b111100000;
				8'b1101101: c <= 9'b1001001;
				8'b100011: c <= 9'b1001010;
				8'b1110101: c <= 9'b10000010;
				8'b1111101: c <= 9'b111101111;
				8'b101001: c <= 9'b110011;
				8'b1010010: c <= 9'b111010000;
				8'b1011000: c <= 9'b11111001;
				8'b101110: c <= 9'b101000100;
				8'b1000001: c <= 9'b110110111;
				default: c <= 9'b0;
			endcase
			9'b1010010 : case(di)
				8'b1000011: c <= 9'b11111;
				8'b101000: c <= 9'b11001100;
				8'b111010: c <= 9'b101000;
				8'b110110: c <= 9'b10000101;
				8'b1100100: c <= 9'b10110101;
				8'b1000000: c <= 9'b11101011;
				8'b1110110: c <= 9'b111100011;
				8'b100101: c <= 9'b100011101;
				8'b101111: c <= 9'b110001011;
				8'b100110: c <= 9'b11100100;
				8'b1100011: c <= 9'b10110100;
				8'b1001000: c <= 9'b111000010;
				8'b111000: c <= 9'b100010000;
				8'b110001: c <= 9'b110010001;
				8'b1010111: c <= 9'b11001;
				8'b1001110: c <= 9'b111100000;
				8'b1101010: c <= 9'b10100;
				8'b1001001: c <= 9'b101011001;
				8'b1100000: c <= 9'b100000110;
				8'b110111: c <= 9'b100000100;
				8'b1011101: c <= 9'b110010110;
				8'b1011011: c <= 9'b1011010;
				8'b111001: c <= 9'b100000010;
				8'b1001010: c <= 9'b111011;
				8'b110011: c <= 9'b1110100;
				8'b1101100: c <= 9'b10011011;
				8'b1110111: c <= 9'b110100101;
				8'b101011: c <= 9'b100000110;
				8'b1101011: c <= 9'b110111;
				8'b111100: c <= 9'b1110010;
				8'b1000111: c <= 9'b101011010;
				8'b1011111: c <= 9'b100111101;
				8'b1110100: c <= 9'b111001111;
				8'b101101: c <= 9'b111001010;
				8'b1010011: c <= 9'b100000101;
				8'b1100001: c <= 9'b111000000;
				8'b110101: c <= 9'b110010100;
				8'b1000100: c <= 9'b111010110;
				8'b1010001: c <= 9'b100000111;
				8'b1010100: c <= 9'b111010000;
				8'b1100110: c <= 9'b10101001;
				8'b101010: c <= 9'b110011010;
				8'b1011110: c <= 9'b111011011;
				8'b1100111: c <= 9'b111110011;
				8'b1011010: c <= 9'b111110011;
				8'b1000010: c <= 9'b111100000;
				8'b111101: c <= 9'b10110001;
				8'b110000: c <= 9'b111000111;
				8'b111110: c <= 9'b100110100;
				8'b1100010: c <= 9'b111111001;
				8'b1110000: c <= 9'b100010110;
				8'b1101001: c <= 9'b111001101;
				8'b1110011: c <= 9'b1110010;
				8'b1001100: c <= 9'b10111001;
				8'b100001: c <= 9'b100001;
				8'b1000110: c <= 9'b111001;
				8'b1110010: c <= 9'b10100010;
				8'b1010000: c <= 9'b100010011;
				8'b1111010: c <= 9'b101010011;
				8'b1010101: c <= 9'b110110111;
				8'b111011: c <= 9'b100100001;
				8'b1001101: c <= 9'b10011011;
				8'b111111: c <= 9'b11100101;
				8'b1101110: c <= 9'b111101010;
				8'b1111011: c <= 9'b11111011;
				8'b1001011: c <= 9'b11111000;
				8'b1101111: c <= 9'b100110;
				8'b1101000: c <= 9'b10001011;
				8'b101100: c <= 9'b110011;
				8'b100100: c <= 9'b110010010;
				8'b1111000: c <= 9'b11110011;
				8'b1000101: c <= 9'b100011101;
				8'b1011001: c <= 9'b10010000;
				8'b110100: c <= 9'b1100100;
				8'b1111001: c <= 9'b101110;
				8'b1110001: c <= 9'b110111110;
				8'b1001111: c <= 9'b1100101;
				8'b1100101: c <= 9'b10011;
				8'b1111110: c <= 9'b101100110;
				8'b1111100: c <= 9'b110110111;
				8'b1010110: c <= 9'b110000101;
				8'b110010: c <= 9'b11100000;
				8'b1101101: c <= 9'b110001111;
				8'b100011: c <= 9'b10001111;
				8'b1110101: c <= 9'b1001;
				8'b1111101: c <= 9'b100001110;
				8'b101001: c <= 9'b1011111;
				8'b1010010: c <= 9'b101100111;
				8'b1011000: c <= 9'b100000010;
				8'b101110: c <= 9'b100001001;
				8'b1000001: c <= 9'b101101010;
				default: c <= 9'b0;
			endcase
			9'b101101011 : case(di)
				8'b1000011: c <= 9'b11101101;
				8'b101000: c <= 9'b110010110;
				8'b111010: c <= 9'b110001011;
				8'b110110: c <= 9'b11111100;
				8'b1100100: c <= 9'b110010001;
				8'b1000000: c <= 9'b100101000;
				8'b1110110: c <= 9'b1011000;
				8'b100101: c <= 9'b10111011;
				8'b101111: c <= 9'b111001111;
				8'b100110: c <= 9'b111111110;
				8'b1100011: c <= 9'b11111101;
				8'b1001000: c <= 9'b111101000;
				8'b111000: c <= 9'b1110000;
				8'b110001: c <= 9'b110010101;
				8'b1010111: c <= 9'b11000100;
				8'b1001110: c <= 9'b100;
				8'b1101010: c <= 9'b1111101;
				8'b1001001: c <= 9'b11101111;
				8'b1100000: c <= 9'b100;
				8'b110111: c <= 9'b10111100;
				8'b1011101: c <= 9'b11110110;
				8'b1011011: c <= 9'b10101111;
				8'b111001: c <= 9'b11100011;
				8'b1001010: c <= 9'b110111010;
				8'b110011: c <= 9'b110001000;
				8'b1101100: c <= 9'b1010000;
				8'b1110111: c <= 9'b10110011;
				8'b101011: c <= 9'b100001100;
				8'b1101011: c <= 9'b110011001;
				8'b111100: c <= 9'b1010000;
				8'b1000111: c <= 9'b1001;
				8'b1011111: c <= 9'b10110;
				8'b1110100: c <= 9'b100110101;
				8'b101101: c <= 9'b10111110;
				8'b1010011: c <= 9'b1000111;
				8'b1100001: c <= 9'b110000111;
				8'b110101: c <= 9'b110010110;
				8'b1000100: c <= 9'b101000011;
				8'b1010001: c <= 9'b11101001;
				8'b1010100: c <= 9'b1001100;
				8'b1100110: c <= 9'b110011001;
				8'b101010: c <= 9'b11100;
				8'b1011110: c <= 9'b110001001;
				8'b1100111: c <= 9'b101110000;
				8'b1011010: c <= 9'b10001001;
				8'b1000010: c <= 9'b100110101;
				8'b111101: c <= 9'b101100101;
				8'b110000: c <= 9'b1100000;
				8'b111110: c <= 9'b10001101;
				8'b1100010: c <= 9'b10110;
				8'b1110000: c <= 9'b10000011;
				8'b1101001: c <= 9'b111011100;
				8'b1110011: c <= 9'b11000000;
				8'b1001100: c <= 9'b10101101;
				8'b100001: c <= 9'b101100001;
				8'b1000110: c <= 9'b110100001;
				8'b1110010: c <= 9'b11111010;
				8'b1010000: c <= 9'b1100010;
				8'b1111010: c <= 9'b101101;
				8'b1010101: c <= 9'b110001001;
				8'b111011: c <= 9'b11111100;
				8'b1001101: c <= 9'b110000111;
				8'b111111: c <= 9'b11110000;
				8'b1101110: c <= 9'b111001010;
				8'b1111011: c <= 9'b100000001;
				8'b1001011: c <= 9'b101111110;
				8'b1101111: c <= 9'b100110010;
				8'b1101000: c <= 9'b11100011;
				8'b101100: c <= 9'b111011101;
				8'b100100: c <= 9'b11001000;
				8'b1111000: c <= 9'b1100011;
				8'b1000101: c <= 9'b110100;
				8'b1011001: c <= 9'b11101001;
				8'b110100: c <= 9'b110101011;
				8'b1111001: c <= 9'b10111100;
				8'b1110001: c <= 9'b111100;
				8'b1001111: c <= 9'b11000011;
				8'b1100101: c <= 9'b11111000;
				8'b1111110: c <= 9'b101011101;
				8'b1111100: c <= 9'b101001;
				8'b1010110: c <= 9'b1011100;
				8'b110010: c <= 9'b110110110;
				8'b1101101: c <= 9'b101100101;
				8'b100011: c <= 9'b1101100;
				8'b1110101: c <= 9'b10111011;
				8'b1111101: c <= 9'b100110;
				8'b101001: c <= 9'b100111110;
				8'b1010010: c <= 9'b1000111;
				8'b1011000: c <= 9'b110001010;
				8'b101110: c <= 9'b100101111;
				8'b1000001: c <= 9'b10000;
				default: c <= 9'b0;
			endcase
			9'b11110000 : case(di)
				8'b1000011: c <= 9'b100100010;
				8'b101000: c <= 9'b101101111;
				8'b111010: c <= 9'b101010110;
				8'b110110: c <= 9'b10001111;
				8'b1100100: c <= 9'b100111;
				8'b1000000: c <= 9'b100010110;
				8'b1110110: c <= 9'b11110110;
				8'b100101: c <= 9'b111011;
				8'b101111: c <= 9'b110110;
				8'b100110: c <= 9'b100010010;
				8'b1100011: c <= 9'b101101110;
				8'b1001000: c <= 9'b11101;
				8'b111000: c <= 9'b110001010;
				8'b110001: c <= 9'b1100110;
				8'b1010111: c <= 9'b10100010;
				8'b1001110: c <= 9'b101011000;
				8'b1101010: c <= 9'b101010101;
				8'b1001001: c <= 9'b111111010;
				8'b1100000: c <= 9'b101011011;
				8'b110111: c <= 9'b101001001;
				8'b1011101: c <= 9'b110000011;
				8'b1011011: c <= 9'b110001101;
				8'b111001: c <= 9'b10111010;
				8'b1001010: c <= 9'b1110100;
				8'b110011: c <= 9'b111010000;
				8'b1101100: c <= 9'b111000100;
				8'b1110111: c <= 9'b1101111;
				8'b101011: c <= 9'b101100110;
				8'b1101011: c <= 9'b110000110;
				8'b111100: c <= 9'b100001011;
				8'b1000111: c <= 9'b1110000;
				8'b1011111: c <= 9'b11100001;
				8'b1110100: c <= 9'b101101110;
				8'b101101: c <= 9'b101100101;
				8'b1010011: c <= 9'b10100011;
				8'b1100001: c <= 9'b11110101;
				8'b110101: c <= 9'b100011101;
				8'b1000100: c <= 9'b1100011;
				8'b1010001: c <= 9'b101111110;
				8'b1010100: c <= 9'b10001010;
				8'b1100110: c <= 9'b1100011;
				8'b101010: c <= 9'b111111;
				8'b1011110: c <= 9'b111001001;
				8'b1100111: c <= 9'b111000010;
				8'b1011010: c <= 9'b100;
				8'b1000010: c <= 9'b110011010;
				8'b111101: c <= 9'b1101001;
				8'b110000: c <= 9'b100101001;
				8'b111110: c <= 9'b110011110;
				8'b1100010: c <= 9'b10101001;
				8'b1110000: c <= 9'b101101110;
				8'b1101001: c <= 9'b1011100;
				8'b1110011: c <= 9'b11000111;
				8'b1001100: c <= 9'b110100000;
				8'b100001: c <= 9'b11111011;
				8'b1000110: c <= 9'b100111101;
				8'b1110010: c <= 9'b101111111;
				8'b1010000: c <= 9'b101001011;
				8'b1111010: c <= 9'b110;
				8'b1010101: c <= 9'b111011100;
				8'b111011: c <= 9'b100110101;
				8'b1001101: c <= 9'b101011010;
				8'b111111: c <= 9'b11101111;
				8'b1101110: c <= 9'b101011001;
				8'b1111011: c <= 9'b1111;
				8'b1001011: c <= 9'b111010100;
				8'b1101111: c <= 9'b110010111;
				8'b1101000: c <= 9'b10000011;
				8'b101100: c <= 9'b11101111;
				8'b100100: c <= 9'b10010;
				8'b1111000: c <= 9'b111010010;
				8'b1000101: c <= 9'b11101;
				8'b1011001: c <= 9'b11011011;
				8'b110100: c <= 9'b101000100;
				8'b1111001: c <= 9'b101101011;
				8'b1110001: c <= 9'b101100;
				8'b1001111: c <= 9'b10001001;
				8'b1100101: c <= 9'b1100101;
				8'b1111110: c <= 9'b100010100;
				8'b1111100: c <= 9'b101100101;
				8'b1010110: c <= 9'b100101111;
				8'b110010: c <= 9'b110101;
				8'b1101101: c <= 9'b110011110;
				8'b100011: c <= 9'b11011110;
				8'b1110101: c <= 9'b101010011;
				8'b1111101: c <= 9'b11010111;
				8'b101001: c <= 9'b1010101;
				8'b1010010: c <= 9'b10001101;
				8'b1011000: c <= 9'b11100011;
				8'b101110: c <= 9'b111010110;
				8'b1000001: c <= 9'b101100101;
				default: c <= 9'b0;
			endcase
			9'b100111101 : case(di)
				8'b1000011: c <= 9'b10101111;
				8'b101000: c <= 9'b11001011;
				8'b111010: c <= 9'b101011000;
				8'b110110: c <= 9'b100110011;
				8'b1100100: c <= 9'b10010100;
				8'b1000000: c <= 9'b11110111;
				8'b1110110: c <= 9'b110110;
				8'b100101: c <= 9'b1010010;
				8'b101111: c <= 9'b100100101;
				8'b100110: c <= 9'b111101010;
				8'b1100011: c <= 9'b10100011;
				8'b1001000: c <= 9'b100111000;
				8'b111000: c <= 9'b11111101;
				8'b110001: c <= 9'b110010110;
				8'b1010111: c <= 9'b101011001;
				8'b1001110: c <= 9'b1011001;
				8'b1101010: c <= 9'b100011000;
				8'b1001001: c <= 9'b11111001;
				8'b1100000: c <= 9'b11000001;
				8'b110111: c <= 9'b10001000;
				8'b1011101: c <= 9'b1100000;
				8'b1011011: c <= 9'b10100010;
				8'b111001: c <= 9'b1000101;
				8'b1001010: c <= 9'b100101001;
				8'b110011: c <= 9'b100000111;
				8'b1101100: c <= 9'b1110011;
				8'b1110111: c <= 9'b1000010;
				8'b101011: c <= 9'b101101100;
				8'b1101011: c <= 9'b10110110;
				8'b111100: c <= 9'b100110100;
				8'b1000111: c <= 9'b110110;
				8'b1011111: c <= 9'b111011001;
				8'b1110100: c <= 9'b1;
				8'b101101: c <= 9'b10000110;
				8'b1010011: c <= 9'b111111110;
				8'b1100001: c <= 9'b10100110;
				8'b110101: c <= 9'b100000101;
				8'b1000100: c <= 9'b10110011;
				8'b1010001: c <= 9'b100001101;
				8'b1010100: c <= 9'b111011100;
				8'b1100110: c <= 9'b11011000;
				8'b101010: c <= 9'b11001010;
				8'b1011110: c <= 9'b1000;
				8'b1100111: c <= 9'b100011011;
				8'b1011010: c <= 9'b111111011;
				8'b1000010: c <= 9'b110111000;
				8'b111101: c <= 9'b10100110;
				8'b110000: c <= 9'b100000011;
				8'b111110: c <= 9'b110111011;
				8'b1100010: c <= 9'b11011010;
				8'b1110000: c <= 9'b11100;
				8'b1101001: c <= 9'b110001100;
				8'b1110011: c <= 9'b110001;
				8'b1001100: c <= 9'b111100001;
				8'b100001: c <= 9'b111100101;
				8'b1000110: c <= 9'b10010011;
				8'b1110010: c <= 9'b1101;
				8'b1010000: c <= 9'b110000001;
				8'b1111010: c <= 9'b11101000;
				8'b1010101: c <= 9'b101110110;
				8'b111011: c <= 9'b1110010;
				8'b1001101: c <= 9'b101100100;
				8'b111111: c <= 9'b1100110;
				8'b1101110: c <= 9'b11001010;
				8'b1111011: c <= 9'b101001100;
				8'b1001011: c <= 9'b10000001;
				8'b1101111: c <= 9'b10100011;
				8'b1101000: c <= 9'b1010010;
				8'b101100: c <= 9'b111011110;
				8'b100100: c <= 9'b110111000;
				8'b1111000: c <= 9'b110010100;
				8'b1000101: c <= 9'b10011001;
				8'b1011001: c <= 9'b11101;
				8'b110100: c <= 9'b10010000;
				8'b1111001: c <= 9'b111111;
				8'b1110001: c <= 9'b101000111;
				8'b1001111: c <= 9'b101011000;
				8'b1100101: c <= 9'b10111010;
				8'b1111110: c <= 9'b100110110;
				8'b1111100: c <= 9'b100001011;
				8'b1010110: c <= 9'b11110010;
				8'b110010: c <= 9'b11010100;
				8'b1101101: c <= 9'b111111111;
				8'b100011: c <= 9'b110001000;
				8'b1110101: c <= 9'b10110110;
				8'b1111101: c <= 9'b110111100;
				8'b101001: c <= 9'b1100000;
				8'b1010010: c <= 9'b100110000;
				8'b1011000: c <= 9'b11011011;
				8'b101110: c <= 9'b10011;
				8'b1000001: c <= 9'b101010101;
				default: c <= 9'b0;
			endcase
			9'b111000000 : case(di)
				8'b1000011: c <= 9'b100100101;
				8'b101000: c <= 9'b101111010;
				8'b111010: c <= 9'b1001000;
				8'b110110: c <= 9'b110011111;
				8'b1100100: c <= 9'b10110101;
				8'b1000000: c <= 9'b11100000;
				8'b1110110: c <= 9'b100000010;
				8'b100101: c <= 9'b100001010;
				8'b101111: c <= 9'b111010111;
				8'b100110: c <= 9'b10000011;
				8'b1100011: c <= 9'b101111110;
				8'b1001000: c <= 9'b111101010;
				8'b111000: c <= 9'b110100010;
				8'b110001: c <= 9'b111111111;
				8'b1010111: c <= 9'b101011110;
				8'b1001110: c <= 9'b10011100;
				8'b1101010: c <= 9'b110010001;
				8'b1001001: c <= 9'b100010100;
				8'b1100000: c <= 9'b100111001;
				8'b110111: c <= 9'b101;
				8'b1011101: c <= 9'b101101011;
				8'b1011011: c <= 9'b110011;
				8'b111001: c <= 9'b100111111;
				8'b1001010: c <= 9'b100101100;
				8'b110011: c <= 9'b110111;
				8'b1101100: c <= 9'b1110101;
				8'b1110111: c <= 9'b100101010;
				8'b101011: c <= 9'b101111110;
				8'b1101011: c <= 9'b11001110;
				8'b111100: c <= 9'b101;
				8'b1000111: c <= 9'b110;
				8'b1011111: c <= 9'b110110110;
				8'b1110100: c <= 9'b101100;
				8'b101101: c <= 9'b11000111;
				8'b1010011: c <= 9'b100111;
				8'b1100001: c <= 9'b10011100;
				8'b110101: c <= 9'b1111011;
				8'b1000100: c <= 9'b100101000;
				8'b1010001: c <= 9'b100011001;
				8'b1010100: c <= 9'b1101001;
				8'b1100110: c <= 9'b11000110;
				8'b101010: c <= 9'b110000110;
				8'b1011110: c <= 9'b101010101;
				8'b1100111: c <= 9'b110011100;
				8'b1011010: c <= 9'b110011100;
				8'b1000010: c <= 9'b101001100;
				8'b111101: c <= 9'b1110111;
				8'b110000: c <= 9'b100110111;
				8'b111110: c <= 9'b100000111;
				8'b1100010: c <= 9'b1100100;
				8'b1110000: c <= 9'b110100111;
				8'b1101001: c <= 9'b111010001;
				8'b1110011: c <= 9'b10111111;
				8'b1001100: c <= 9'b101010101;
				8'b100001: c <= 9'b10101001;
				8'b1000110: c <= 9'b111011111;
				8'b1110010: c <= 9'b11110000;
				8'b1010000: c <= 9'b111111110;
				8'b1111010: c <= 9'b110111011;
				8'b1010101: c <= 9'b1111101;
				8'b111011: c <= 9'b110011110;
				8'b1001101: c <= 9'b100111101;
				8'b111111: c <= 9'b1100010;
				8'b1101110: c <= 9'b111010001;
				8'b1111011: c <= 9'b100111011;
				8'b1001011: c <= 9'b1010011;
				8'b1101111: c <= 9'b100101101;
				8'b1101000: c <= 9'b101;
				8'b101100: c <= 9'b110001001;
				8'b100100: c <= 9'b10101001;
				8'b1111000: c <= 9'b110000;
				8'b1000101: c <= 9'b11100000;
				8'b1011001: c <= 9'b110010111;
				8'b110100: c <= 9'b111000101;
				8'b1111001: c <= 9'b10010100;
				8'b1110001: c <= 9'b100110101;
				8'b1001111: c <= 9'b100101011;
				8'b1100101: c <= 9'b11000000;
				8'b1111110: c <= 9'b10101100;
				8'b1111100: c <= 9'b100011000;
				8'b1010110: c <= 9'b100000011;
				8'b110010: c <= 9'b111111101;
				8'b1101101: c <= 9'b110100101;
				8'b100011: c <= 9'b1011000;
				8'b1110101: c <= 9'b1001100;
				8'b1111101: c <= 9'b100010010;
				8'b101001: c <= 9'b11001111;
				8'b1010010: c <= 9'b1111011;
				8'b1011000: c <= 9'b10001000;
				8'b101110: c <= 9'b110110111;
				8'b1000001: c <= 9'b100010010;
				default: c <= 9'b0;
			endcase
			9'b10111011 : case(di)
				8'b1000011: c <= 9'b1010110;
				8'b101000: c <= 9'b101110010;
				8'b111010: c <= 9'b11110001;
				8'b110110: c <= 9'b1111010;
				8'b1100100: c <= 9'b100110100;
				8'b1000000: c <= 9'b101101111;
				8'b1110110: c <= 9'b110101101;
				8'b100101: c <= 9'b111100001;
				8'b101111: c <= 9'b11000000;
				8'b100110: c <= 9'b111111;
				8'b1100011: c <= 9'b111111110;
				8'b1001000: c <= 9'b10010100;
				8'b111000: c <= 9'b110011010;
				8'b110001: c <= 9'b100000110;
				8'b1010111: c <= 9'b110111011;
				8'b1001110: c <= 9'b10010001;
				8'b1101010: c <= 9'b11111101;
				8'b1001001: c <= 9'b10001110;
				8'b1100000: c <= 9'b1100001;
				8'b110111: c <= 9'b100110100;
				8'b1011101: c <= 9'b101001010;
				8'b1011011: c <= 9'b11010010;
				8'b111001: c <= 9'b110100011;
				8'b1001010: c <= 9'b110111001;
				8'b110011: c <= 9'b11111100;
				8'b1101100: c <= 9'b1100110;
				8'b1110111: c <= 9'b111011111;
				8'b101011: c <= 9'b1111111;
				8'b1101011: c <= 9'b11010101;
				8'b111100: c <= 9'b11100101;
				8'b1000111: c <= 9'b1011;
				8'b1011111: c <= 9'b11110101;
				8'b1110100: c <= 9'b10010001;
				8'b101101: c <= 9'b101001011;
				8'b1010011: c <= 9'b11000100;
				8'b1100001: c <= 9'b11111;
				8'b110101: c <= 9'b1011001;
				8'b1000100: c <= 9'b111110011;
				8'b1010001: c <= 9'b111100001;
				8'b1010100: c <= 9'b10011100;
				8'b1100110: c <= 9'b10100;
				8'b101010: c <= 9'b110000111;
				8'b1011110: c <= 9'b111100110;
				8'b1100111: c <= 9'b111100011;
				8'b1011010: c <= 9'b10101111;
				8'b1000010: c <= 9'b1000011;
				8'b111101: c <= 9'b100001011;
				8'b110000: c <= 9'b101100111;
				8'b111110: c <= 9'b110101100;
				8'b1100010: c <= 9'b10101011;
				8'b1110000: c <= 9'b111111001;
				8'b1101001: c <= 9'b11100000;
				8'b1110011: c <= 9'b11010100;
				8'b1001100: c <= 9'b1001011;
				8'b100001: c <= 9'b10000010;
				8'b1000110: c <= 9'b110100010;
				8'b1110010: c <= 9'b11110100;
				8'b1010000: c <= 9'b11101000;
				8'b1111010: c <= 9'b101101110;
				8'b1010101: c <= 9'b11100;
				8'b111011: c <= 9'b110111110;
				8'b1001101: c <= 9'b100010110;
				8'b111111: c <= 9'b111101101;
				8'b1101110: c <= 9'b1001001;
				8'b1111011: c <= 9'b11011011;
				8'b1001011: c <= 9'b1011000;
				8'b1101111: c <= 9'b111111000;
				8'b1101000: c <= 9'b10011101;
				8'b101100: c <= 9'b10000000;
				8'b100100: c <= 9'b11000011;
				8'b1111000: c <= 9'b101111001;
				8'b1000101: c <= 9'b11101;
				8'b1011001: c <= 9'b11101011;
				8'b110100: c <= 9'b1000010;
				8'b1111001: c <= 9'b110111111;
				8'b1110001: c <= 9'b10010011;
				8'b1001111: c <= 9'b111011010;
				8'b1100101: c <= 9'b101110010;
				8'b1111110: c <= 9'b111111000;
				8'b1111100: c <= 9'b111110000;
				8'b1010110: c <= 9'b110010001;
				8'b110010: c <= 9'b1101111;
				8'b1101101: c <= 9'b100000101;
				8'b100011: c <= 9'b1010000;
				8'b1110101: c <= 9'b1110101;
				8'b1111101: c <= 9'b10110001;
				8'b101001: c <= 9'b1000110;
				8'b1010010: c <= 9'b11010101;
				8'b1011000: c <= 9'b111011010;
				8'b101110: c <= 9'b101;
				8'b1000001: c <= 9'b1010001;
				default: c <= 9'b0;
			endcase
			9'b11001110 : case(di)
				8'b1000011: c <= 9'b10000111;
				8'b101000: c <= 9'b111100001;
				8'b111010: c <= 9'b110010001;
				8'b110110: c <= 9'b100110100;
				8'b1100100: c <= 9'b1011010;
				8'b1000000: c <= 9'b101001;
				8'b1110110: c <= 9'b101100100;
				8'b100101: c <= 9'b11100001;
				8'b101111: c <= 9'b11100101;
				8'b100110: c <= 9'b1000011;
				8'b1100011: c <= 9'b111111011;
				8'b1001000: c <= 9'b111110011;
				8'b111000: c <= 9'b110001110;
				8'b110001: c <= 9'b11111101;
				8'b1010111: c <= 9'b1011010;
				8'b1001110: c <= 9'b1101100;
				8'b1101010: c <= 9'b111110001;
				8'b1001001: c <= 9'b100111011;
				8'b1100000: c <= 9'b11010011;
				8'b110111: c <= 9'b101011101;
				8'b1011101: c <= 9'b101011110;
				8'b1011011: c <= 9'b100001001;
				8'b111001: c <= 9'b101101101;
				8'b1001010: c <= 9'b11110111;
				8'b110011: c <= 9'b10011111;
				8'b1101100: c <= 9'b110011011;
				8'b1110111: c <= 9'b1111111;
				8'b101011: c <= 9'b100101010;
				8'b1101011: c <= 9'b1100;
				8'b111100: c <= 9'b11100111;
				8'b1000111: c <= 9'b100000101;
				8'b1011111: c <= 9'b11000010;
				8'b1110100: c <= 9'b111101;
				8'b101101: c <= 9'b11011110;
				8'b1010011: c <= 9'b1011001;
				8'b1100001: c <= 9'b110101100;
				8'b110101: c <= 9'b11100;
				8'b1000100: c <= 9'b110101010;
				8'b1010001: c <= 9'b11010100;
				8'b1010100: c <= 9'b111110001;
				8'b1100110: c <= 9'b1011001;
				8'b101010: c <= 9'b110011100;
				8'b1011110: c <= 9'b100111000;
				8'b1100111: c <= 9'b1010111;
				8'b1011010: c <= 9'b11011110;
				8'b1000010: c <= 9'b101110010;
				8'b111101: c <= 9'b11100011;
				8'b110000: c <= 9'b11010111;
				8'b111110: c <= 9'b111010000;
				8'b1100010: c <= 9'b1111100;
				8'b1110000: c <= 9'b100111111;
				8'b1101001: c <= 9'b101100100;
				8'b1110011: c <= 9'b1001011;
				8'b1001100: c <= 9'b110110100;
				8'b100001: c <= 9'b111111101;
				8'b1000110: c <= 9'b110111001;
				8'b1110010: c <= 9'b1001110;
				8'b1010000: c <= 9'b110011111;
				8'b1111010: c <= 9'b100111010;
				8'b1010101: c <= 9'b11000110;
				8'b111011: c <= 9'b1100010;
				8'b1001101: c <= 9'b101101011;
				8'b111111: c <= 9'b110000011;
				8'b1101110: c <= 9'b11101001;
				8'b1111011: c <= 9'b10111011;
				8'b1001011: c <= 9'b10001000;
				8'b1101111: c <= 9'b10101100;
				8'b1101000: c <= 9'b100011101;
				8'b101100: c <= 9'b100110110;
				8'b100100: c <= 9'b11011000;
				8'b1111000: c <= 9'b110100000;
				8'b1000101: c <= 9'b11101011;
				8'b1011001: c <= 9'b10001111;
				8'b110100: c <= 9'b110100;
				8'b1111001: c <= 9'b101010101;
				8'b1110001: c <= 9'b100011111;
				8'b1001111: c <= 9'b100001111;
				8'b1100101: c <= 9'b11001;
				8'b1111110: c <= 9'b11010101;
				8'b1111100: c <= 9'b101011000;
				8'b1010110: c <= 9'b10010101;
				8'b110010: c <= 9'b111011011;
				8'b1101101: c <= 9'b100011001;
				8'b100011: c <= 9'b10111101;
				8'b1110101: c <= 9'b1111110;
				8'b1111101: c <= 9'b11100010;
				8'b101001: c <= 9'b110000;
				8'b1010010: c <= 9'b111010001;
				8'b1011000: c <= 9'b1;
				8'b101110: c <= 9'b11111100;
				8'b1000001: c <= 9'b1100101;
				default: c <= 9'b0;
			endcase
			9'b100001010 : case(di)
				8'b1000011: c <= 9'b111000010;
				8'b101000: c <= 9'b1010001;
				8'b111010: c <= 9'b1000010;
				8'b110110: c <= 9'b10111001;
				8'b1100100: c <= 9'b110010010;
				8'b1000000: c <= 9'b10111110;
				8'b1110110: c <= 9'b11;
				8'b100101: c <= 9'b1010101;
				8'b101111: c <= 9'b10010;
				8'b100110: c <= 9'b1100100;
				8'b1100011: c <= 9'b100101101;
				8'b1001000: c <= 9'b111011001;
				8'b111000: c <= 9'b11001101;
				8'b110001: c <= 9'b1100000;
				8'b1010111: c <= 9'b10011;
				8'b1001110: c <= 9'b111101001;
				8'b1101010: c <= 9'b11110101;
				8'b1001001: c <= 9'b101010111;
				8'b1100000: c <= 9'b11111;
				8'b110111: c <= 9'b111101010;
				8'b1011101: c <= 9'b10001010;
				8'b1011011: c <= 9'b100100001;
				8'b111001: c <= 9'b1111;
				8'b1001010: c <= 9'b111001;
				8'b110011: c <= 9'b111001110;
				8'b1101100: c <= 9'b110011101;
				8'b1110111: c <= 9'b111110101;
				8'b101011: c <= 9'b10011010;
				8'b1101011: c <= 9'b100001001;
				8'b111100: c <= 9'b101100001;
				8'b1000111: c <= 9'b111011001;
				8'b1011111: c <= 9'b1011111;
				8'b1110100: c <= 9'b11100011;
				8'b101101: c <= 9'b111000111;
				8'b1010011: c <= 9'b110100001;
				8'b1100001: c <= 9'b110111010;
				8'b110101: c <= 9'b111010000;
				8'b1000100: c <= 9'b10001110;
				8'b1010001: c <= 9'b11010010;
				8'b1010100: c <= 9'b100010011;
				8'b1100110: c <= 9'b101101010;
				8'b101010: c <= 9'b101010110;
				8'b1011110: c <= 9'b100010111;
				8'b1100111: c <= 9'b101011110;
				8'b1011010: c <= 9'b1111001;
				8'b1000010: c <= 9'b11101000;
				8'b111101: c <= 9'b110101001;
				8'b110000: c <= 9'b100010100;
				8'b111110: c <= 9'b111100100;
				8'b1100010: c <= 9'b100111110;
				8'b1110000: c <= 9'b11110111;
				8'b1101001: c <= 9'b11111000;
				8'b1110011: c <= 9'b101100001;
				8'b1001100: c <= 9'b1100010;
				8'b100001: c <= 9'b100100001;
				8'b1000110: c <= 9'b100101001;
				8'b1110010: c <= 9'b11110100;
				8'b1010000: c <= 9'b100100000;
				8'b1111010: c <= 9'b11101;
				8'b1010101: c <= 9'b1001111;
				8'b111011: c <= 9'b11111100;
				8'b1001101: c <= 9'b100100;
				8'b111111: c <= 9'b10101110;
				8'b1101110: c <= 9'b10101100;
				8'b1111011: c <= 9'b111001111;
				8'b1001011: c <= 9'b10101011;
				8'b1101111: c <= 9'b10110001;
				8'b1101000: c <= 9'b10000111;
				8'b101100: c <= 9'b1100000;
				8'b100100: c <= 9'b10011001;
				8'b1111000: c <= 9'b100100110;
				8'b1000101: c <= 9'b111010100;
				8'b1011001: c <= 9'b101010001;
				8'b110100: c <= 9'b10111;
				8'b1111001: c <= 9'b100001101;
				8'b1110001: c <= 9'b111100010;
				8'b1001111: c <= 9'b110001010;
				8'b1100101: c <= 9'b11000110;
				8'b1111110: c <= 9'b1101001;
				8'b1111100: c <= 9'b100001010;
				8'b1010110: c <= 9'b1011010;
				8'b110010: c <= 9'b1101111;
				8'b1101101: c <= 9'b1110010;
				8'b100011: c <= 9'b10000101;
				8'b1110101: c <= 9'b11;
				8'b1111101: c <= 9'b10010;
				8'b101001: c <= 9'b100101001;
				8'b1010010: c <= 9'b1111011;
				8'b1011000: c <= 9'b11101101;
				8'b101110: c <= 9'b111100;
				8'b1000001: c <= 9'b110010011;
				default: c <= 9'b0;
			endcase
			9'b100011000 : case(di)
				8'b1000011: c <= 9'b100110100;
				8'b101000: c <= 9'b1111101;
				8'b111010: c <= 9'b101010001;
				8'b110110: c <= 9'b111000;
				8'b1100100: c <= 9'b110110111;
				8'b1000000: c <= 9'b1011110;
				8'b1110110: c <= 9'b1111;
				8'b100101: c <= 9'b1111101;
				8'b101111: c <= 9'b110001011;
				8'b100110: c <= 9'b100100000;
				8'b1100011: c <= 9'b10010000;
				8'b1001000: c <= 9'b100111001;
				8'b111000: c <= 9'b1100100;
				8'b110001: c <= 9'b110101110;
				8'b1010111: c <= 9'b100100111;
				8'b1001110: c <= 9'b101110100;
				8'b1101010: c <= 9'b100101101;
				8'b1001001: c <= 9'b110101101;
				8'b1100000: c <= 9'b110010010;
				8'b110111: c <= 9'b111001111;
				8'b1011101: c <= 9'b111100000;
				8'b1011011: c <= 9'b100001101;
				8'b111001: c <= 9'b11011001;
				8'b1001010: c <= 9'b10000111;
				8'b110011: c <= 9'b100101010;
				8'b1101100: c <= 9'b111010110;
				8'b1110111: c <= 9'b100110;
				8'b101011: c <= 9'b101000011;
				8'b1101011: c <= 9'b111111000;
				8'b111100: c <= 9'b100010010;
				8'b1000111: c <= 9'b110010111;
				8'b1011111: c <= 9'b111011100;
				8'b1110100: c <= 9'b10110110;
				8'b101101: c <= 9'b111011011;
				8'b1010011: c <= 9'b10001110;
				8'b1100001: c <= 9'b110110110;
				8'b110101: c <= 9'b110100010;
				8'b1000100: c <= 9'b100010110;
				8'b1010001: c <= 9'b110010011;
				8'b1010100: c <= 9'b10000;
				8'b1100110: c <= 9'b111101010;
				8'b101010: c <= 9'b101101001;
				8'b1011110: c <= 9'b11010000;
				8'b1100111: c <= 9'b10011111;
				8'b1011010: c <= 9'b101011000;
				8'b1000010: c <= 9'b101111110;
				8'b111101: c <= 9'b10001011;
				8'b110000: c <= 9'b111011001;
				8'b111110: c <= 9'b10011;
				8'b1100010: c <= 9'b11111000;
				8'b1110000: c <= 9'b100110;
				8'b1101001: c <= 9'b100100111;
				8'b1110011: c <= 9'b1110011;
				8'b1001100: c <= 9'b110101011;
				8'b100001: c <= 9'b10011;
				8'b1000110: c <= 9'b1000001;
				8'b1110010: c <= 9'b11101011;
				8'b1010000: c <= 9'b10100010;
				8'b1111010: c <= 9'b10010001;
				8'b1010101: c <= 9'b101011;
				8'b111011: c <= 9'b1111000;
				8'b1001101: c <= 9'b10111000;
				8'b111111: c <= 9'b110100000;
				8'b1101110: c <= 9'b100001110;
				8'b1111011: c <= 9'b1110000;
				8'b1001011: c <= 9'b10000111;
				8'b1101111: c <= 9'b110101;
				8'b1101000: c <= 9'b100111010;
				8'b101100: c <= 9'b11010010;
				8'b100100: c <= 9'b11010011;
				8'b1111000: c <= 9'b101001000;
				8'b1000101: c <= 9'b11110101;
				8'b1011001: c <= 9'b10111111;
				8'b110100: c <= 9'b101100001;
				8'b1111001: c <= 9'b110111110;
				8'b1110001: c <= 9'b10111101;
				8'b1001111: c <= 9'b110110000;
				8'b1100101: c <= 9'b101101110;
				8'b1111110: c <= 9'b100101100;
				8'b1111100: c <= 9'b110011101;
				8'b1010110: c <= 9'b100111010;
				8'b110010: c <= 9'b101010100;
				8'b1101101: c <= 9'b111000010;
				8'b100011: c <= 9'b100101010;
				8'b1110101: c <= 9'b110111;
				8'b1111101: c <= 9'b10011000;
				8'b101001: c <= 9'b100000100;
				8'b1010010: c <= 9'b100010000;
				8'b1011000: c <= 9'b100001110;
				8'b101110: c <= 9'b100011111;
				8'b1000001: c <= 9'b101011110;
				default: c <= 9'b0;
			endcase
			9'b11111101 : case(di)
				8'b1000011: c <= 9'b1111;
				8'b101000: c <= 9'b110111010;
				8'b111010: c <= 9'b11101111;
				8'b110110: c <= 9'b110110110;
				8'b1100100: c <= 9'b1100010;
				8'b1000000: c <= 9'b101000101;
				8'b1110110: c <= 9'b1100101;
				8'b100101: c <= 9'b110101101;
				8'b101111: c <= 9'b100101101;
				8'b100110: c <= 9'b111100001;
				8'b1100011: c <= 9'b111101010;
				8'b1001000: c <= 9'b11000010;
				8'b111000: c <= 9'b10111;
				8'b110001: c <= 9'b110111110;
				8'b1010111: c <= 9'b11110011;
				8'b1001110: c <= 9'b10101;
				8'b1101010: c <= 9'b111111000;
				8'b1001001: c <= 9'b110000;
				8'b1100000: c <= 9'b1001010;
				8'b110111: c <= 9'b1010110;
				8'b1011101: c <= 9'b100000110;
				8'b1011011: c <= 9'b101101110;
				8'b111001: c <= 9'b111001001;
				8'b1001010: c <= 9'b11101001;
				8'b110011: c <= 9'b10011010;
				8'b1101100: c <= 9'b11011100;
				8'b1110111: c <= 9'b110;
				8'b101011: c <= 9'b111000010;
				8'b1101011: c <= 9'b101010101;
				8'b111100: c <= 9'b1110010;
				8'b1000111: c <= 9'b101011001;
				8'b1011111: c <= 9'b10111100;
				8'b1110100: c <= 9'b10001101;
				8'b101101: c <= 9'b101111010;
				8'b1010011: c <= 9'b100100010;
				8'b1100001: c <= 9'b1001010;
				8'b110101: c <= 9'b110101111;
				8'b1000100: c <= 9'b100010000;
				8'b1010001: c <= 9'b100000101;
				8'b1010100: c <= 9'b10000111;
				8'b1100110: c <= 9'b100111110;
				8'b101010: c <= 9'b100111101;
				8'b1011110: c <= 9'b11101000;
				8'b1100111: c <= 9'b10000101;
				8'b1011010: c <= 9'b110010011;
				8'b1000010: c <= 9'b10011011;
				8'b111101: c <= 9'b111100010;
				8'b110000: c <= 9'b10000111;
				8'b111110: c <= 9'b1101110;
				8'b1100010: c <= 9'b11100100;
				8'b1110000: c <= 9'b11100;
				8'b1101001: c <= 9'b110010010;
				8'b1110011: c <= 9'b101111111;
				8'b1001100: c <= 9'b11100011;
				8'b100001: c <= 9'b110010;
				8'b1000110: c <= 9'b11001101;
				8'b1110010: c <= 9'b101011001;
				8'b1010000: c <= 9'b111110110;
				8'b1111010: c <= 9'b100;
				8'b1010101: c <= 9'b111100001;
				8'b111011: c <= 9'b11100110;
				8'b1001101: c <= 9'b1001;
				8'b111111: c <= 9'b10000010;
				8'b1101110: c <= 9'b110111100;
				8'b1111011: c <= 9'b110011010;
				8'b1001011: c <= 9'b11110001;
				8'b1101111: c <= 9'b11110011;
				8'b1101000: c <= 9'b111010100;
				8'b101100: c <= 9'b101000010;
				8'b100100: c <= 9'b1111100;
				8'b1111000: c <= 9'b10011000;
				8'b1000101: c <= 9'b11001111;
				8'b1011001: c <= 9'b11101011;
				8'b110100: c <= 9'b100111001;
				8'b1111001: c <= 9'b10111110;
				8'b1110001: c <= 9'b110100101;
				8'b1001111: c <= 9'b100011001;
				8'b1100101: c <= 9'b11110001;
				8'b1111110: c <= 9'b111111101;
				8'b1111100: c <= 9'b1001001;
				8'b1010110: c <= 9'b1010111;
				8'b110010: c <= 9'b10011100;
				8'b1101101: c <= 9'b1110001;
				8'b100011: c <= 9'b1101010;
				8'b1110101: c <= 9'b101101011;
				8'b1111101: c <= 9'b100100001;
				8'b101001: c <= 9'b101011001;
				8'b1010010: c <= 9'b10101011;
				8'b1011000: c <= 9'b101110100;
				8'b101110: c <= 9'b111011101;
				8'b1000001: c <= 9'b1000001;
				default: c <= 9'b0;
			endcase
			9'b11100110 : case(di)
				8'b1000011: c <= 9'b101101001;
				8'b101000: c <= 9'b110011010;
				8'b111010: c <= 9'b101101010;
				8'b110110: c <= 9'b10110110;
				8'b1100100: c <= 9'b110000010;
				8'b1000000: c <= 9'b101101100;
				8'b1110110: c <= 9'b110100111;
				8'b100101: c <= 9'b11100100;
				8'b101111: c <= 9'b101101010;
				8'b100110: c <= 9'b110010010;
				8'b1100011: c <= 9'b100110110;
				8'b1001000: c <= 9'b111111101;
				8'b111000: c <= 9'b10100011;
				8'b110001: c <= 9'b100010000;
				8'b1010111: c <= 9'b1010011;
				8'b1001110: c <= 9'b11110000;
				8'b1101010: c <= 9'b110111111;
				8'b1001001: c <= 9'b11010100;
				8'b1100000: c <= 9'b101100010;
				8'b110111: c <= 9'b11111001;
				8'b1011101: c <= 9'b110;
				8'b1011011: c <= 9'b10110011;
				8'b111001: c <= 9'b110100100;
				8'b1001010: c <= 9'b10;
				8'b110011: c <= 9'b101010;
				8'b1101100: c <= 9'b110001101;
				8'b1110111: c <= 9'b11110111;
				8'b101011: c <= 9'b110000101;
				8'b1101011: c <= 9'b101100101;
				8'b111100: c <= 9'b111001101;
				8'b1000111: c <= 9'b111101101;
				8'b1011111: c <= 9'b110000000;
				8'b1110100: c <= 9'b110000000;
				8'b101101: c <= 9'b110110;
				8'b1010011: c <= 9'b110010001;
				8'b1100001: c <= 9'b111100111;
				8'b110101: c <= 9'b111110110;
				8'b1000100: c <= 9'b101111000;
				8'b1010001: c <= 9'b110001;
				8'b1010100: c <= 9'b1100100;
				8'b1100110: c <= 9'b101011000;
				8'b101010: c <= 9'b10110100;
				8'b1011110: c <= 9'b101001111;
				8'b1100111: c <= 9'b100011000;
				8'b1011010: c <= 9'b101000110;
				8'b1000010: c <= 9'b10000;
				8'b111101: c <= 9'b111110001;
				8'b110000: c <= 9'b111100100;
				8'b111110: c <= 9'b11000111;
				8'b1100010: c <= 9'b110111001;
				8'b1110000: c <= 9'b111011001;
				8'b1101001: c <= 9'b110001001;
				8'b1110011: c <= 9'b11111;
				8'b1001100: c <= 9'b1111101;
				8'b100001: c <= 9'b110011100;
				8'b1000110: c <= 9'b1111001;
				8'b1110010: c <= 9'b11010101;
				8'b1010000: c <= 9'b101110000;
				8'b1111010: c <= 9'b11010010;
				8'b1010101: c <= 9'b110111010;
				8'b111011: c <= 9'b111001110;
				8'b1001101: c <= 9'b11011000;
				8'b111111: c <= 9'b101101110;
				8'b1101110: c <= 9'b1011100;
				8'b1111011: c <= 9'b110100;
				8'b1001011: c <= 9'b10011;
				8'b1101111: c <= 9'b11100001;
				8'b1101000: c <= 9'b101000;
				8'b101100: c <= 9'b101101011;
				8'b100100: c <= 9'b1111;
				8'b1111000: c <= 9'b111000000;
				8'b1000101: c <= 9'b1011000;
				8'b1011001: c <= 9'b11100001;
				8'b110100: c <= 9'b100000000;
				8'b1111001: c <= 9'b11111101;
				8'b1110001: c <= 9'b10110;
				8'b1001111: c <= 9'b101111001;
				8'b1100101: c <= 9'b111001101;
				8'b1111110: c <= 9'b110010110;
				8'b1111100: c <= 9'b110100111;
				8'b1010110: c <= 9'b110000110;
				8'b110010: c <= 9'b11001000;
				8'b1101101: c <= 9'b100011000;
				8'b100011: c <= 9'b1;
				8'b1110101: c <= 9'b101011110;
				8'b1111101: c <= 9'b110010;
				8'b101001: c <= 9'b11100110;
				8'b1010010: c <= 9'b100010010;
				8'b1011000: c <= 9'b10011011;
				8'b101110: c <= 9'b111101100;
				8'b1000001: c <= 9'b100011000;
				default: c <= 9'b0;
			endcase
			9'b111100001 : case(di)
				8'b1000011: c <= 9'b100010;
				8'b101000: c <= 9'b1100101;
				8'b111010: c <= 9'b100111000;
				8'b110110: c <= 9'b10010;
				8'b1100100: c <= 9'b110001001;
				8'b1000000: c <= 9'b101101001;
				8'b1110110: c <= 9'b111000010;
				8'b100101: c <= 9'b100111101;
				8'b101111: c <= 9'b101111110;
				8'b100110: c <= 9'b100010;
				8'b1100011: c <= 9'b110100111;
				8'b1001000: c <= 9'b10001011;
				8'b111000: c <= 9'b101101000;
				8'b110001: c <= 9'b110001110;
				8'b1010111: c <= 9'b110000010;
				8'b1001110: c <= 9'b1100001;
				8'b1101010: c <= 9'b111001100;
				8'b1001001: c <= 9'b111110110;
				8'b1100000: c <= 9'b10100011;
				8'b110111: c <= 9'b11010001;
				8'b1011101: c <= 9'b10001100;
				8'b1011011: c <= 9'b1101101;
				8'b111001: c <= 9'b100100;
				8'b1001010: c <= 9'b111100111;
				8'b110011: c <= 9'b101100011;
				8'b1101100: c <= 9'b100111010;
				8'b1110111: c <= 9'b1110111;
				8'b101011: c <= 9'b100010;
				8'b1101011: c <= 9'b100010010;
				8'b111100: c <= 9'b1000010;
				8'b1000111: c <= 9'b11100011;
				8'b1011111: c <= 9'b1100000;
				8'b1110100: c <= 9'b111000111;
				8'b101101: c <= 9'b111111;
				8'b1010011: c <= 9'b10;
				8'b1100001: c <= 9'b1011111;
				8'b110101: c <= 9'b110010001;
				8'b1000100: c <= 9'b1111;
				8'b1010001: c <= 9'b1110100;
				8'b1010100: c <= 9'b10101101;
				8'b1100110: c <= 9'b100100001;
				8'b101010: c <= 9'b111001001;
				8'b1011110: c <= 9'b100100001;
				8'b1100111: c <= 9'b11011000;
				8'b1011010: c <= 9'b111011101;
				8'b1000010: c <= 9'b1111100;
				8'b111101: c <= 9'b100000000;
				8'b110000: c <= 9'b111010111;
				8'b111110: c <= 9'b100111000;
				8'b1100010: c <= 9'b1101001;
				8'b1110000: c <= 9'b100110;
				8'b1101001: c <= 9'b1001000;
				8'b1110011: c <= 9'b111000;
				8'b1001100: c <= 9'b110110;
				8'b100001: c <= 9'b10110;
				8'b1000110: c <= 9'b100101111;
				8'b1110010: c <= 9'b111;
				8'b1010000: c <= 9'b1111001;
				8'b1111010: c <= 9'b100000001;
				8'b1010101: c <= 9'b11101001;
				8'b111011: c <= 9'b111100001;
				8'b1001101: c <= 9'b1001110;
				8'b111111: c <= 9'b111001011;
				8'b1101110: c <= 9'b100;
				8'b1111011: c <= 9'b100000101;
				8'b1001011: c <= 9'b101000111;
				8'b1101111: c <= 9'b1001110;
				8'b1101000: c <= 9'b11011000;
				8'b101100: c <= 9'b110101100;
				8'b100100: c <= 9'b1010101;
				8'b1111000: c <= 9'b100100000;
				8'b1000101: c <= 9'b111101010;
				8'b1011001: c <= 9'b101100101;
				8'b110100: c <= 9'b101000;
				8'b1111001: c <= 9'b1000011;
				8'b1110001: c <= 9'b1111100;
				8'b1001111: c <= 9'b111100001;
				8'b1100101: c <= 9'b10111101;
				8'b1111110: c <= 9'b10111011;
				8'b1111100: c <= 9'b1010111;
				8'b1010110: c <= 9'b10111011;
				8'b110010: c <= 9'b111000;
				8'b1101101: c <= 9'b111101100;
				8'b100011: c <= 9'b10111010;
				8'b1110101: c <= 9'b110001100;
				8'b1111101: c <= 9'b100100000;
				8'b101001: c <= 9'b11110000;
				8'b1010010: c <= 9'b101000010;
				8'b1011000: c <= 9'b111111111;
				8'b101110: c <= 9'b1100010;
				8'b1000001: c <= 9'b101111010;
				default: c <= 9'b0;
			endcase
			9'b1010011 : case(di)
				8'b1000011: c <= 9'b110100101;
				8'b101000: c <= 9'b10011111;
				8'b111010: c <= 9'b110001011;
				8'b110110: c <= 9'b110111111;
				8'b1100100: c <= 9'b10101000;
				8'b1000000: c <= 9'b11001110;
				8'b1110110: c <= 9'b100111111;
				8'b100101: c <= 9'b10101;
				8'b101111: c <= 9'b110011;
				8'b100110: c <= 9'b111111;
				8'b1100011: c <= 9'b101100;
				8'b1001000: c <= 9'b100001;
				8'b111000: c <= 9'b11110111;
				8'b110001: c <= 9'b1010101;
				8'b1010111: c <= 9'b101001110;
				8'b1001110: c <= 9'b111111000;
				8'b1101010: c <= 9'b11100011;
				8'b1001001: c <= 9'b101101010;
				8'b1100000: c <= 9'b11000000;
				8'b110111: c <= 9'b100110100;
				8'b1011101: c <= 9'b111000100;
				8'b1011011: c <= 9'b100000010;
				8'b111001: c <= 9'b101110010;
				8'b1001010: c <= 9'b100111110;
				8'b110011: c <= 9'b110000001;
				8'b1101100: c <= 9'b111111011;
				8'b1110111: c <= 9'b1100111;
				8'b101011: c <= 9'b10100101;
				8'b1101011: c <= 9'b110010110;
				8'b111100: c <= 9'b10100110;
				8'b1000111: c <= 9'b111010;
				8'b1011111: c <= 9'b10010101;
				8'b1110100: c <= 9'b100000111;
				8'b101101: c <= 9'b11111101;
				8'b1010011: c <= 9'b101100101;
				8'b1100001: c <= 9'b110001100;
				8'b110101: c <= 9'b1000010;
				8'b1000100: c <= 9'b100111011;
				8'b1010001: c <= 9'b11110001;
				8'b1010100: c <= 9'b110101111;
				8'b1100110: c <= 9'b110010110;
				8'b101010: c <= 9'b111011011;
				8'b1011110: c <= 9'b10111011;
				8'b1100111: c <= 9'b100101010;
				8'b1011010: c <= 9'b100110;
				8'b1000010: c <= 9'b110001;
				8'b111101: c <= 9'b10001100;
				8'b110000: c <= 9'b11101011;
				8'b111110: c <= 9'b11111010;
				8'b1100010: c <= 9'b1010001;
				8'b1110000: c <= 9'b101101010;
				8'b1101001: c <= 9'b10110101;
				8'b1110011: c <= 9'b101110001;
				8'b1001100: c <= 9'b10101110;
				8'b100001: c <= 9'b11011000;
				8'b1000110: c <= 9'b11110001;
				8'b1110010: c <= 9'b100001110;
				8'b1010000: c <= 9'b1011100;
				8'b1111010: c <= 9'b110110000;
				8'b1010101: c <= 9'b111100;
				8'b111011: c <= 9'b11110011;
				8'b1001101: c <= 9'b11100101;
				8'b111111: c <= 9'b11000011;
				8'b1101110: c <= 9'b110001010;
				8'b1111011: c <= 9'b11000;
				8'b1001011: c <= 9'b11000111;
				8'b1101111: c <= 9'b11100111;
				8'b1101000: c <= 9'b100101000;
				8'b101100: c <= 9'b111100000;
				8'b100100: c <= 9'b100000100;
				8'b1111000: c <= 9'b1000011;
				8'b1000101: c <= 9'b10010111;
				8'b1011001: c <= 9'b1110;
				8'b110100: c <= 9'b101000011;
				8'b1111001: c <= 9'b110110011;
				8'b1110001: c <= 9'b1010010;
				8'b1001111: c <= 9'b11011;
				8'b1100101: c <= 9'b110100011;
				8'b1111110: c <= 9'b101010;
				8'b1111100: c <= 9'b101010111;
				8'b1010110: c <= 9'b10101111;
				8'b110010: c <= 9'b10000111;
				8'b1101101: c <= 9'b100011000;
				8'b100011: c <= 9'b1001010;
				8'b1110101: c <= 9'b101111110;
				8'b1111101: c <= 9'b111000011;
				8'b101001: c <= 9'b1101010;
				8'b1010010: c <= 9'b1001111;
				8'b1011000: c <= 9'b10001001;
				8'b101110: c <= 9'b110110110;
				8'b1000001: c <= 9'b100111101;
				default: c <= 9'b0;
			endcase
			9'b1101 : case(di)
				8'b1000011: c <= 9'b101100110;
				8'b101000: c <= 9'b10000001;
				8'b111010: c <= 9'b101001001;
				8'b110110: c <= 9'b1001011;
				8'b1100100: c <= 9'b101110111;
				8'b1000000: c <= 9'b111011010;
				8'b1110110: c <= 9'b111011101;
				8'b100101: c <= 9'b110010010;
				8'b101111: c <= 9'b110111110;
				8'b100110: c <= 9'b111001110;
				8'b1100011: c <= 9'b110011010;
				8'b1001000: c <= 9'b100011;
				8'b111000: c <= 9'b101110;
				8'b110001: c <= 9'b1101001;
				8'b1010111: c <= 9'b111000111;
				8'b1001110: c <= 9'b100001;
				8'b1101010: c <= 9'b1101110;
				8'b1001001: c <= 9'b11111010;
				8'b1100000: c <= 9'b101000011;
				8'b110111: c <= 9'b111001;
				8'b1011101: c <= 9'b100110010;
				8'b1011011: c <= 9'b100111001;
				8'b111001: c <= 9'b101110110;
				8'b1001010: c <= 9'b111010100;
				8'b110011: c <= 9'b10011;
				8'b1101100: c <= 9'b11110100;
				8'b1110111: c <= 9'b100001001;
				8'b101011: c <= 9'b10001100;
				8'b1101011: c <= 9'b11001110;
				8'b111100: c <= 9'b11101011;
				8'b1000111: c <= 9'b10111101;
				8'b1011111: c <= 9'b1101110;
				8'b1110100: c <= 9'b1010001;
				8'b101101: c <= 9'b110101100;
				8'b1010011: c <= 9'b111101001;
				8'b1100001: c <= 9'b110011011;
				8'b110101: c <= 9'b100111;
				8'b1000100: c <= 9'b11111;
				8'b1010001: c <= 9'b111100;
				8'b1010100: c <= 9'b11110;
				8'b1100110: c <= 9'b101001000;
				8'b101010: c <= 9'b110000011;
				8'b1011110: c <= 9'b10110010;
				8'b1100111: c <= 9'b100100110;
				8'b1011010: c <= 9'b111101111;
				8'b1000010: c <= 9'b11001110;
				8'b111101: c <= 9'b110100100;
				8'b110000: c <= 9'b1100101;
				8'b111110: c <= 9'b110111000;
				8'b1100010: c <= 9'b10001111;
				8'b1110000: c <= 9'b100000010;
				8'b1101001: c <= 9'b10010100;
				8'b1110011: c <= 9'b11111101;
				8'b1001100: c <= 9'b111000101;
				8'b100001: c <= 9'b101110001;
				8'b1000110: c <= 9'b10010100;
				8'b1110010: c <= 9'b101100100;
				8'b1010000: c <= 9'b10110;
				8'b1111010: c <= 9'b11010010;
				8'b1010101: c <= 9'b100010101;
				8'b111011: c <= 9'b100001;
				8'b1001101: c <= 9'b11111101;
				8'b111111: c <= 9'b111011011;
				8'b1101110: c <= 9'b1000000;
				8'b1111011: c <= 9'b100011001;
				8'b1001011: c <= 9'b1111000;
				8'b1101111: c <= 9'b100111000;
				8'b1101000: c <= 9'b110100;
				8'b101100: c <= 9'b111010001;
				8'b100100: c <= 9'b111101101;
				8'b1111000: c <= 9'b110111010;
				8'b1000101: c <= 9'b11101000;
				8'b1011001: c <= 9'b11010;
				8'b110100: c <= 9'b10110100;
				8'b1111001: c <= 9'b10000001;
				8'b1110001: c <= 9'b100000111;
				8'b1001111: c <= 9'b111011110;
				8'b1100101: c <= 9'b110111001;
				8'b1111110: c <= 9'b110011001;
				8'b1111100: c <= 9'b111010000;
				8'b1010110: c <= 9'b111000010;
				8'b110010: c <= 9'b111000111;
				8'b1101101: c <= 9'b110001;
				8'b100011: c <= 9'b10110101;
				8'b1110101: c <= 9'b11010111;
				8'b1111101: c <= 9'b111101100;
				8'b101001: c <= 9'b1100000;
				8'b1010010: c <= 9'b110111011;
				8'b1011000: c <= 9'b110101001;
				8'b101110: c <= 9'b100101101;
				8'b1000001: c <= 9'b10010111;
				default: c <= 9'b0;
			endcase
			9'b1100001 : case(di)
				8'b1000011: c <= 9'b111100101;
				8'b101000: c <= 9'b1;
				8'b111010: c <= 9'b100011010;
				8'b110110: c <= 9'b11111101;
				8'b1100100: c <= 9'b101001001;
				8'b1000000: c <= 9'b101001100;
				8'b1110110: c <= 9'b100111001;
				8'b100101: c <= 9'b10000001;
				8'b101111: c <= 9'b10001001;
				8'b100110: c <= 9'b110011111;
				8'b1100011: c <= 9'b100000001;
				8'b1001000: c <= 9'b1110;
				8'b111000: c <= 9'b100110101;
				8'b110001: c <= 9'b10010110;
				8'b1010111: c <= 9'b11110011;
				8'b1001110: c <= 9'b10110001;
				8'b1101010: c <= 9'b111011110;
				8'b1001001: c <= 9'b101111010;
				8'b1100000: c <= 9'b1001;
				8'b110111: c <= 9'b1010001;
				8'b1011101: c <= 9'b1011;
				8'b1011011: c <= 9'b10001111;
				8'b111001: c <= 9'b1001;
				8'b1001010: c <= 9'b110101110;
				8'b110011: c <= 9'b1001000;
				8'b1101100: c <= 9'b110010100;
				8'b1110111: c <= 9'b101011111;
				8'b101011: c <= 9'b111100110;
				8'b1101011: c <= 9'b11000010;
				8'b111100: c <= 9'b111001;
				8'b1000111: c <= 9'b100110000;
				8'b1011111: c <= 9'b1000110;
				8'b1110100: c <= 9'b1000000;
				8'b101101: c <= 9'b101001001;
				8'b1010011: c <= 9'b101001001;
				8'b1100001: c <= 9'b100001110;
				8'b110101: c <= 9'b101101001;
				8'b1000100: c <= 9'b10111100;
				8'b1010001: c <= 9'b100100000;
				8'b1010100: c <= 9'b111011111;
				8'b1100110: c <= 9'b101001110;
				8'b101010: c <= 9'b10010011;
				8'b1011110: c <= 9'b11110110;
				8'b1100111: c <= 9'b100111111;
				8'b1011010: c <= 9'b111000000;
				8'b1000010: c <= 9'b110011;
				8'b111101: c <= 9'b10000110;
				8'b110000: c <= 9'b110011001;
				8'b111110: c <= 9'b100100011;
				8'b1100010: c <= 9'b100110111;
				8'b1110000: c <= 9'b100000100;
				8'b1101001: c <= 9'b111100101;
				8'b1110011: c <= 9'b1101010;
				8'b1001100: c <= 9'b101100110;
				8'b100001: c <= 9'b111100111;
				8'b1000110: c <= 9'b1011110;
				8'b1110010: c <= 9'b110100100;
				8'b1010000: c <= 9'b110101010;
				8'b1111010: c <= 9'b100100111;
				8'b1010101: c <= 9'b110101001;
				8'b111011: c <= 9'b11111000;
				8'b1001101: c <= 9'b110101100;
				8'b111111: c <= 9'b111010111;
				8'b1101110: c <= 9'b1111000;
				8'b1111011: c <= 9'b111001111;
				8'b1001011: c <= 9'b10011111;
				8'b1101111: c <= 9'b10011001;
				8'b1101000: c <= 9'b100110100;
				8'b101100: c <= 9'b1;
				8'b100100: c <= 9'b1010011;
				8'b1111000: c <= 9'b110111011;
				8'b1000101: c <= 9'b101011010;
				8'b1011001: c <= 9'b111000010;
				8'b110100: c <= 9'b101000011;
				8'b1111001: c <= 9'b10010011;
				8'b1110001: c <= 9'b10011010;
				8'b1001111: c <= 9'b10000101;
				8'b1100101: c <= 9'b101011001;
				8'b1111110: c <= 9'b111001101;
				8'b1111100: c <= 9'b110111;
				8'b1010110: c <= 9'b100001101;
				8'b110010: c <= 9'b1000001;
				8'b1101101: c <= 9'b10001100;
				8'b100011: c <= 9'b110001111;
				8'b1110101: c <= 9'b10011011;
				8'b1111101: c <= 9'b100010110;
				8'b101001: c <= 9'b111010111;
				8'b1010010: c <= 9'b11110;
				8'b1011000: c <= 9'b101001001;
				8'b101110: c <= 9'b100101101;
				8'b1000001: c <= 9'b110100001;
				default: c <= 9'b0;
			endcase
			9'b10001111 : case(di)
				8'b1000011: c <= 9'b110011000;
				8'b101000: c <= 9'b111000100;
				8'b111010: c <= 9'b111011110;
				8'b110110: c <= 9'b11010100;
				8'b1100100: c <= 9'b101110010;
				8'b1000000: c <= 9'b10110011;
				8'b1110110: c <= 9'b101010111;
				8'b100101: c <= 9'b111100111;
				8'b101111: c <= 9'b100101011;
				8'b100110: c <= 9'b1101100;
				8'b1100011: c <= 9'b11110000;
				8'b1001000: c <= 9'b11100111;
				8'b111000: c <= 9'b101100;
				8'b110001: c <= 9'b10010101;
				8'b1010111: c <= 9'b100111000;
				8'b1001110: c <= 9'b100011111;
				8'b1101010: c <= 9'b111111110;
				8'b1001001: c <= 9'b11100011;
				8'b1100000: c <= 9'b101011;
				8'b110111: c <= 9'b111111011;
				8'b1011101: c <= 9'b11110011;
				8'b1011011: c <= 9'b101010001;
				8'b111001: c <= 9'b11001101;
				8'b1001010: c <= 9'b1001000;
				8'b110011: c <= 9'b110110110;
				8'b1101100: c <= 9'b110010110;
				8'b1110111: c <= 9'b110111010;
				8'b101011: c <= 9'b100011010;
				8'b1101011: c <= 9'b11110100;
				8'b111100: c <= 9'b10;
				8'b1000111: c <= 9'b111101111;
				8'b1011111: c <= 9'b101101001;
				8'b1110100: c <= 9'b110011011;
				8'b101101: c <= 9'b11001000;
				8'b1010011: c <= 9'b1110000;
				8'b1100001: c <= 9'b111101110;
				8'b110101: c <= 9'b111100100;
				8'b1000100: c <= 9'b100101110;
				8'b1010001: c <= 9'b110101011;
				8'b1010100: c <= 9'b11101011;
				8'b1100110: c <= 9'b110011101;
				8'b101010: c <= 9'b101100110;
				8'b1011110: c <= 9'b1001101;
				8'b1100111: c <= 9'b111100001;
				8'b1011010: c <= 9'b111001110;
				8'b1000010: c <= 9'b111100011;
				8'b111101: c <= 9'b101101001;
				8'b110000: c <= 9'b100000111;
				8'b111110: c <= 9'b101000111;
				8'b1100010: c <= 9'b101011111;
				8'b1110000: c <= 9'b111000111;
				8'b1101001: c <= 9'b100101;
				8'b1110011: c <= 9'b100100000;
				8'b1001100: c <= 9'b11011001;
				8'b100001: c <= 9'b10101000;
				8'b1000110: c <= 9'b11;
				8'b1110010: c <= 9'b1110001;
				8'b1010000: c <= 9'b110010001;
				8'b1111010: c <= 9'b11011001;
				8'b1010101: c <= 9'b11111010;
				8'b111011: c <= 9'b11110111;
				8'b1001101: c <= 9'b1011100;
				8'b111111: c <= 9'b10100111;
				8'b1101110: c <= 9'b11000100;
				8'b1111011: c <= 9'b111001001;
				8'b1001011: c <= 9'b101111110;
				8'b1101111: c <= 9'b10010;
				8'b1101000: c <= 9'b1100100;
				8'b101100: c <= 9'b11011101;
				8'b100100: c <= 9'b100000110;
				8'b1111000: c <= 9'b101;
				8'b1000101: c <= 9'b11100;
				8'b1011001: c <= 9'b110111100;
				8'b110100: c <= 9'b100100001;
				8'b1111001: c <= 9'b11101;
				8'b1110001: c <= 9'b1100111;
				8'b1001111: c <= 9'b10101111;
				8'b1100101: c <= 9'b1101101;
				8'b1111110: c <= 9'b101101;
				8'b1111100: c <= 9'b110101101;
				8'b1010110: c <= 9'b110001;
				8'b110010: c <= 9'b10110010;
				8'b1101101: c <= 9'b1110001;
				8'b100011: c <= 9'b100010011;
				8'b1110101: c <= 9'b110111010;
				8'b1111101: c <= 9'b11110101;
				8'b101001: c <= 9'b100110011;
				8'b1010010: c <= 9'b100110101;
				8'b1011000: c <= 9'b11000010;
				8'b101110: c <= 9'b101001100;
				8'b1000001: c <= 9'b111001010;
				default: c <= 9'b0;
			endcase
			9'b111000011 : case(di)
				8'b1000011: c <= 9'b10011001;
				8'b101000: c <= 9'b101001001;
				8'b111010: c <= 9'b10011010;
				8'b110110: c <= 9'b110100010;
				8'b1100100: c <= 9'b100111010;
				8'b1000000: c <= 9'b110101;
				8'b1110110: c <= 9'b111000111;
				8'b100101: c <= 9'b111000;
				8'b101111: c <= 9'b11010011;
				8'b100110: c <= 9'b1000;
				8'b1100011: c <= 9'b11010000;
				8'b1001000: c <= 9'b100011001;
				8'b111000: c <= 9'b10000001;
				8'b110001: c <= 9'b1010001;
				8'b1010111: c <= 9'b110000000;
				8'b1001110: c <= 9'b111000100;
				8'b1101010: c <= 9'b110111;
				8'b1001001: c <= 9'b110100000;
				8'b1100000: c <= 9'b110000000;
				8'b110111: c <= 9'b101111001;
				8'b1011101: c <= 9'b100010;
				8'b1011011: c <= 9'b111000011;
				8'b111001: c <= 9'b11110000;
				8'b1001010: c <= 9'b1101101;
				8'b110011: c <= 9'b101100010;
				8'b1101100: c <= 9'b100111101;
				8'b1110111: c <= 9'b111101100;
				8'b101011: c <= 9'b1101001;
				8'b1101011: c <= 9'b111010111;
				8'b111100: c <= 9'b111111000;
				8'b1000111: c <= 9'b111011110;
				8'b1011111: c <= 9'b11111010;
				8'b1110100: c <= 9'b111011011;
				8'b101101: c <= 9'b101001010;
				8'b1010011: c <= 9'b110001011;
				8'b1100001: c <= 9'b11101011;
				8'b110101: c <= 9'b100011001;
				8'b1000100: c <= 9'b10101011;
				8'b1010001: c <= 9'b10101100;
				8'b1010100: c <= 9'b101011001;
				8'b1100110: c <= 9'b100010;
				8'b101010: c <= 9'b100000010;
				8'b1011110: c <= 9'b110000110;
				8'b1100111: c <= 9'b101001100;
				8'b1011010: c <= 9'b110011001;
				8'b1000010: c <= 9'b110110111;
				8'b111101: c <= 9'b11111001;
				8'b110000: c <= 9'b111100001;
				8'b111110: c <= 9'b10001000;
				8'b1100010: c <= 9'b101100101;
				8'b1110000: c <= 9'b10101111;
				8'b1101001: c <= 9'b110001100;
				8'b1110011: c <= 9'b101000101;
				8'b1001100: c <= 9'b101010110;
				8'b100001: c <= 9'b1011111;
				8'b1000110: c <= 9'b100101101;
				8'b1110010: c <= 9'b101011000;
				8'b1010000: c <= 9'b101101101;
				8'b1111010: c <= 9'b1000111;
				8'b1010101: c <= 9'b100100;
				8'b111011: c <= 9'b110010101;
				8'b1001101: c <= 9'b101000100;
				8'b111111: c <= 9'b110011101;
				8'b1101110: c <= 9'b10111011;
				8'b1111011: c <= 9'b11001010;
				8'b1001011: c <= 9'b1010111;
				8'b1101111: c <= 9'b1110101;
				8'b1101000: c <= 9'b111010110;
				8'b101100: c <= 9'b101111010;
				8'b100100: c <= 9'b110101100;
				8'b1111000: c <= 9'b101100110;
				8'b1000101: c <= 9'b1011100;
				8'b1011001: c <= 9'b10010101;
				8'b110100: c <= 9'b11011000;
				8'b1111001: c <= 9'b100011010;
				8'b1110001: c <= 9'b110000001;
				8'b1001111: c <= 9'b10101101;
				8'b1100101: c <= 9'b111001001;
				8'b1111110: c <= 9'b11101000;
				8'b1111100: c <= 9'b11;
				8'b1010110: c <= 9'b1101010;
				8'b110010: c <= 9'b100011101;
				8'b1101101: c <= 9'b110000010;
				8'b100011: c <= 9'b1011;
				8'b1110101: c <= 9'b1101;
				8'b1111101: c <= 9'b11000110;
				8'b101001: c <= 9'b11001000;
				8'b1010010: c <= 9'b101100010;
				8'b1011000: c <= 9'b110000011;
				8'b101110: c <= 9'b11100;
				8'b1000001: c <= 9'b110001;
				default: c <= 9'b0;
			endcase
			9'b101111010 : case(di)
				8'b1000011: c <= 9'b110011100;
				8'b101000: c <= 9'b11001101;
				8'b111010: c <= 9'b10010111;
				8'b110110: c <= 9'b11001110;
				8'b1100100: c <= 9'b10100101;
				8'b1000000: c <= 9'b100110010;
				8'b1110110: c <= 9'b11111101;
				8'b100101: c <= 9'b10101111;
				8'b101111: c <= 9'b100110011;
				8'b100110: c <= 9'b11000;
				8'b1100011: c <= 9'b110111011;
				8'b1001000: c <= 9'b10100000;
				8'b111000: c <= 9'b100;
				8'b110001: c <= 9'b100101001;
				8'b1010111: c <= 9'b1010101;
				8'b1001110: c <= 9'b110011101;
				8'b1101010: c <= 9'b111;
				8'b1001001: c <= 9'b110110011;
				8'b1100000: c <= 9'b10010011;
				8'b110111: c <= 9'b10110001;
				8'b1011101: c <= 9'b1111000;
				8'b1011011: c <= 9'b110101011;
				8'b111001: c <= 9'b10000000;
				8'b1001010: c <= 9'b10100;
				8'b110011: c <= 9'b1101111;
				8'b1101100: c <= 9'b110110010;
				8'b1110111: c <= 9'b101101;
				8'b101011: c <= 9'b111000010;
				8'b1101011: c <= 9'b111011010;
				8'b111100: c <= 9'b101011101;
				8'b1000111: c <= 9'b10011001;
				8'b1011111: c <= 9'b100110100;
				8'b1110100: c <= 9'b111100100;
				8'b101101: c <= 9'b100100011;
				8'b1010011: c <= 9'b10010;
				8'b1100001: c <= 9'b10010;
				8'b110101: c <= 9'b110101100;
				8'b1000100: c <= 9'b11000100;
				8'b1010001: c <= 9'b1101111;
				8'b1010100: c <= 9'b11011110;
				8'b1100110: c <= 9'b11001111;
				8'b101010: c <= 9'b110110100;
				8'b1011110: c <= 9'b11011;
				8'b1100111: c <= 9'b100010;
				8'b1011010: c <= 9'b111001110;
				8'b1000010: c <= 9'b10110;
				8'b111101: c <= 9'b111010110;
				8'b110000: c <= 9'b100111000;
				8'b111110: c <= 9'b101110000;
				8'b1100010: c <= 9'b11011;
				8'b1110000: c <= 9'b111010110;
				8'b1101001: c <= 9'b111001100;
				8'b1110011: c <= 9'b111111110;
				8'b1001100: c <= 9'b1001100;
				8'b100001: c <= 9'b11111011;
				8'b1000110: c <= 9'b111010100;
				8'b1110010: c <= 9'b111111111;
				8'b1010000: c <= 9'b11011010;
				8'b1111010: c <= 9'b1100000;
				8'b1010101: c <= 9'b101010;
				8'b111011: c <= 9'b110001000;
				8'b1001101: c <= 9'b111001101;
				8'b111111: c <= 9'b11101000;
				8'b1101110: c <= 9'b100110110;
				8'b1111011: c <= 9'b111001110;
				8'b1001011: c <= 9'b110111111;
				8'b1101111: c <= 9'b1101101;
				8'b1101000: c <= 9'b101010;
				8'b101100: c <= 9'b110111010;
				8'b100100: c <= 9'b10011;
				8'b1111000: c <= 9'b100000011;
				8'b1000101: c <= 9'b10010001;
				8'b1011001: c <= 9'b11110010;
				8'b110100: c <= 9'b11101011;
				8'b1111001: c <= 9'b1100;
				8'b1110001: c <= 9'b1100;
				8'b1001111: c <= 9'b10011001;
				8'b1100101: c <= 9'b10101110;
				8'b1111110: c <= 9'b11111000;
				8'b1111100: c <= 9'b110000010;
				8'b1010110: c <= 9'b111011101;
				8'b110010: c <= 9'b111000101;
				8'b1101101: c <= 9'b100110000;
				8'b100011: c <= 9'b100100;
				8'b1110101: c <= 9'b11011;
				8'b1111101: c <= 9'b1110111;
				8'b101001: c <= 9'b110110100;
				8'b1010010: c <= 9'b1101110;
				8'b1011000: c <= 9'b110111001;
				8'b101110: c <= 9'b11101100;
				8'b1000001: c <= 9'b100001100;
				default: c <= 9'b0;
			endcase
			9'b10001010 : case(di)
				8'b1000011: c <= 9'b100001010;
				8'b101000: c <= 9'b101110100;
				8'b111010: c <= 9'b1101111;
				8'b110110: c <= 9'b101000011;
				8'b1100100: c <= 9'b100101100;
				8'b1000000: c <= 9'b101100000;
				8'b1110110: c <= 9'b111001111;
				8'b100101: c <= 9'b111000011;
				8'b101111: c <= 9'b101101101;
				8'b100110: c <= 9'b11100100;
				8'b1100011: c <= 9'b111000000;
				8'b1001000: c <= 9'b11;
				8'b111000: c <= 9'b110001001;
				8'b110001: c <= 9'b101010100;
				8'b1010111: c <= 9'b10101;
				8'b1001110: c <= 9'b11110011;
				8'b1101010: c <= 9'b110000000;
				8'b1001001: c <= 9'b11010111;
				8'b1100000: c <= 9'b100000011;
				8'b110111: c <= 9'b100101011;
				8'b1011101: c <= 9'b11010111;
				8'b1011011: c <= 9'b10000011;
				8'b111001: c <= 9'b100111001;
				8'b1001010: c <= 9'b100001110;
				8'b110011: c <= 9'b111000;
				8'b1101100: c <= 9'b110001111;
				8'b1110111: c <= 9'b110111000;
				8'b101011: c <= 9'b11001101;
				8'b1101011: c <= 9'b11011010;
				8'b111100: c <= 9'b101011010;
				8'b1000111: c <= 9'b111101101;
				8'b1011111: c <= 9'b11111;
				8'b1110100: c <= 9'b10001010;
				8'b101101: c <= 9'b110011001;
				8'b1010011: c <= 9'b1100001;
				8'b1100001: c <= 9'b10011100;
				8'b110101: c <= 9'b10010101;
				8'b1000100: c <= 9'b11101;
				8'b1010001: c <= 9'b1011001;
				8'b1010100: c <= 9'b100000011;
				8'b1100110: c <= 9'b11110011;
				8'b101010: c <= 9'b1110000;
				8'b1011110: c <= 9'b111010111;
				8'b1100111: c <= 9'b111111101;
				8'b1011010: c <= 9'b111010110;
				8'b1000010: c <= 9'b110100001;
				8'b111101: c <= 9'b110001011;
				8'b110000: c <= 9'b110010111;
				8'b111110: c <= 9'b110101100;
				8'b1100010: c <= 9'b100000110;
				8'b1110000: c <= 9'b11100010;
				8'b1101001: c <= 9'b110111111;
				8'b1110011: c <= 9'b101000001;
				8'b1001100: c <= 9'b100000001;
				8'b100001: c <= 9'b1110111;
				8'b1000110: c <= 9'b10011000;
				8'b1110010: c <= 9'b10111111;
				8'b1010000: c <= 9'b10011001;
				8'b1111010: c <= 9'b110100111;
				8'b1010101: c <= 9'b110101100;
				8'b111011: c <= 9'b1001000;
				8'b1001101: c <= 9'b11101111;
				8'b111111: c <= 9'b100011011;
				8'b1101110: c <= 9'b11;
				8'b1111011: c <= 9'b10010111;
				8'b1001011: c <= 9'b101110110;
				8'b1101111: c <= 9'b111011010;
				8'b1101000: c <= 9'b111001100;
				8'b101100: c <= 9'b111001;
				8'b100100: c <= 9'b10101011;
				8'b1111000: c <= 9'b11111;
				8'b1000101: c <= 9'b111010001;
				8'b1011001: c <= 9'b110010110;
				8'b110100: c <= 9'b11000001;
				8'b1111001: c <= 9'b101001;
				8'b1110001: c <= 9'b1100100;
				8'b1001111: c <= 9'b111010100;
				8'b1100101: c <= 9'b1001111;
				8'b1111110: c <= 9'b1111111;
				8'b1111100: c <= 9'b1110;
				8'b1010110: c <= 9'b110010011;
				8'b110010: c <= 9'b1010101;
				8'b1101101: c <= 9'b101000011;
				8'b100011: c <= 9'b10001110;
				8'b1110101: c <= 9'b101010;
				8'b1111101: c <= 9'b10001100;
				8'b101001: c <= 9'b111101110;
				8'b1010010: c <= 9'b111000011;
				8'b1011000: c <= 9'b110001011;
				8'b101110: c <= 9'b10100111;
				8'b1000001: c <= 9'b100011010;
				default: c <= 9'b0;
			endcase
			9'b1101001 : case(di)
				8'b1000011: c <= 9'b101111000;
				8'b101000: c <= 9'b101001;
				8'b111010: c <= 9'b111010010;
				8'b110110: c <= 9'b1000;
				8'b1100100: c <= 9'b10100011;
				8'b1000000: c <= 9'b11100111;
				8'b1110110: c <= 9'b10001111;
				8'b100101: c <= 9'b101100001;
				8'b101111: c <= 9'b10010111;
				8'b100110: c <= 9'b1111010;
				8'b1100011: c <= 9'b100011111;
				8'b1001000: c <= 9'b11001011;
				8'b111000: c <= 9'b11000;
				8'b110001: c <= 9'b10110101;
				8'b1010111: c <= 9'b101111000;
				8'b1001110: c <= 9'b101100100;
				8'b1101010: c <= 9'b100001010;
				8'b1001001: c <= 9'b101000100;
				8'b1100000: c <= 9'b101000110;
				8'b110111: c <= 9'b110010001;
				8'b1011101: c <= 9'b101101001;
				8'b1011011: c <= 9'b111110011;
				8'b111001: c <= 9'b10110100;
				8'b1001010: c <= 9'b100101000;
				8'b110011: c <= 9'b10110010;
				8'b1101100: c <= 9'b111000011;
				8'b1110111: c <= 9'b110111011;
				8'b101011: c <= 9'b110001111;
				8'b1101011: c <= 9'b110001101;
				8'b111100: c <= 9'b100001110;
				8'b1000111: c <= 9'b110100101;
				8'b1011111: c <= 9'b101100000;
				8'b1110100: c <= 9'b111001111;
				8'b101101: c <= 9'b100110010;
				8'b1010011: c <= 9'b11111101;
				8'b1100001: c <= 9'b1000101;
				8'b110101: c <= 9'b1100111;
				8'b1000100: c <= 9'b11110100;
				8'b1010001: c <= 9'b101000110;
				8'b1010100: c <= 9'b101000010;
				8'b1100110: c <= 9'b10011001;
				8'b101010: c <= 9'b10100110;
				8'b1011110: c <= 9'b10011011;
				8'b1100111: c <= 9'b100001100;
				8'b1011010: c <= 9'b101101101;
				8'b1000010: c <= 9'b101101;
				8'b111101: c <= 9'b110110;
				8'b110000: c <= 9'b100010001;
				8'b111110: c <= 9'b111011100;
				8'b1100010: c <= 9'b101010100;
				8'b1110000: c <= 9'b11011;
				8'b1101001: c <= 9'b10000110;
				8'b1110011: c <= 9'b110011001;
				8'b1001100: c <= 9'b1100101;
				8'b100001: c <= 9'b111011110;
				8'b1000110: c <= 9'b101101110;
				8'b1110010: c <= 9'b1110101;
				8'b1010000: c <= 9'b10000;
				8'b1111010: c <= 9'b101001110;
				8'b1010101: c <= 9'b100101111;
				8'b111011: c <= 9'b100110010;
				8'b1001101: c <= 9'b111011001;
				8'b111111: c <= 9'b110001011;
				8'b1101110: c <= 9'b101011000;
				8'b1111011: c <= 9'b10100011;
				8'b1001011: c <= 9'b11111000;
				8'b1101111: c <= 9'b10100111;
				8'b1101000: c <= 9'b111011011;
				8'b101100: c <= 9'b111001110;
				8'b100100: c <= 9'b10000010;
				8'b1111000: c <= 9'b101001;
				8'b1000101: c <= 9'b100000000;
				8'b1011001: c <= 9'b110000001;
				8'b110100: c <= 9'b10111101;
				8'b1111001: c <= 9'b100110000;
				8'b1110001: c <= 9'b1010011;
				8'b1001111: c <= 9'b11010100;
				8'b1100101: c <= 9'b111011011;
				8'b1111110: c <= 9'b110100;
				8'b1111100: c <= 9'b10001110;
				8'b1010110: c <= 9'b11111010;
				8'b110010: c <= 9'b111111010;
				8'b1101101: c <= 9'b110101;
				8'b100011: c <= 9'b100110010;
				8'b1110101: c <= 9'b110111111;
				8'b1111101: c <= 9'b100000100;
				8'b101001: c <= 9'b11000;
				8'b1010010: c <= 9'b11110101;
				8'b1011000: c <= 9'b10011100;
				8'b101110: c <= 9'b11001011;
				8'b1000001: c <= 9'b11001101;
				default: c <= 9'b0;
			endcase
			9'b10100110 : case(di)
				8'b1000011: c <= 9'b10001110;
				8'b101000: c <= 9'b101000011;
				8'b111010: c <= 9'b1100011;
				8'b110110: c <= 9'b101010001;
				8'b1100100: c <= 9'b100110100;
				8'b1000000: c <= 9'b111110000;
				8'b1110110: c <= 9'b10000111;
				8'b100101: c <= 9'b100011000;
				8'b101111: c <= 9'b11110100;
				8'b100110: c <= 9'b100110101;
				8'b1100011: c <= 9'b101101110;
				8'b1001000: c <= 9'b10011;
				8'b111000: c <= 9'b1110111;
				8'b110001: c <= 9'b100;
				8'b1010111: c <= 9'b101110000;
				8'b1001110: c <= 9'b1000111;
				8'b1101010: c <= 9'b11001101;
				8'b1001001: c <= 9'b11101100;
				8'b1100000: c <= 9'b110010100;
				8'b110111: c <= 9'b11001;
				8'b1011101: c <= 9'b11111010;
				8'b1011011: c <= 9'b111100101;
				8'b111001: c <= 9'b110101100;
				8'b1001010: c <= 9'b10100000;
				8'b110011: c <= 9'b101110010;
				8'b1101100: c <= 9'b101110100;
				8'b1110111: c <= 9'b1111110;
				8'b101011: c <= 9'b1010111;
				8'b1101011: c <= 9'b101101000;
				8'b111100: c <= 9'b100000001;
				8'b1000111: c <= 9'b110000010;
				8'b1011111: c <= 9'b1000001;
				8'b1110100: c <= 9'b1101000;
				8'b101101: c <= 9'b10110010;
				8'b1010011: c <= 9'b10011001;
				8'b1100001: c <= 9'b100101111;
				8'b110101: c <= 9'b101111111;
				8'b1000100: c <= 9'b100111000;
				8'b1010001: c <= 9'b111000010;
				8'b1010100: c <= 9'b110001;
				8'b1100110: c <= 9'b100111;
				8'b101010: c <= 9'b1011110;
				8'b1011110: c <= 9'b110000110;
				8'b1100111: c <= 9'b111000111;
				8'b1011010: c <= 9'b10001010;
				8'b1000010: c <= 9'b10001110;
				8'b111101: c <= 9'b11010010;
				8'b110000: c <= 9'b10000101;
				8'b111110: c <= 9'b101001;
				8'b1100010: c <= 9'b100011;
				8'b1110000: c <= 9'b11;
				8'b1101001: c <= 9'b1010010;
				8'b1110011: c <= 9'b110001000;
				8'b1001100: c <= 9'b11100111;
				8'b100001: c <= 9'b10000011;
				8'b1000110: c <= 9'b101010;
				8'b1110010: c <= 9'b111100;
				8'b1010000: c <= 9'b1001;
				8'b1111010: c <= 9'b1100101;
				8'b1010101: c <= 9'b10111001;
				8'b111011: c <= 9'b1000111;
				8'b1001101: c <= 9'b11000001;
				8'b111111: c <= 9'b1100010;
				8'b1101110: c <= 9'b101011000;
				8'b1111011: c <= 9'b111100000;
				8'b1001011: c <= 9'b1010000;
				8'b1101111: c <= 9'b1011010;
				8'b1101000: c <= 9'b10101101;
				8'b101100: c <= 9'b110010011;
				8'b100100: c <= 9'b110001110;
				8'b1111000: c <= 9'b101101010;
				8'b1000101: c <= 9'b101010100;
				8'b1011001: c <= 9'b110000111;
				8'b110100: c <= 9'b101100100;
				8'b1111001: c <= 9'b101110001;
				8'b1110001: c <= 9'b110001000;
				8'b1001111: c <= 9'b110100110;
				8'b1100101: c <= 9'b100101001;
				8'b1111110: c <= 9'b10100111;
				8'b1111100: c <= 9'b1000010;
				8'b1010110: c <= 9'b10101110;
				8'b110010: c <= 9'b11111;
				8'b1101101: c <= 9'b10110101;
				8'b100011: c <= 9'b1001000;
				8'b1110101: c <= 9'b111110001;
				8'b1111101: c <= 9'b100101101;
				8'b101001: c <= 9'b111100011;
				8'b1010010: c <= 9'b1000111;
				8'b1011000: c <= 9'b11001010;
				8'b101110: c <= 9'b101001100;
				8'b1000001: c <= 9'b100000100;
				default: c <= 9'b0;
			endcase
			9'b110111111 : case(di)
				8'b1000011: c <= 9'b110000;
				8'b101000: c <= 9'b110000000;
				8'b111010: c <= 9'b111000011;
				8'b110110: c <= 9'b101010010;
				8'b1100100: c <= 9'b11000011;
				8'b1000000: c <= 9'b11010;
				8'b1110110: c <= 9'b110101010;
				8'b100101: c <= 9'b101001100;
				8'b101111: c <= 9'b11010000;
				8'b100110: c <= 9'b110111;
				8'b1100011: c <= 9'b1100;
				8'b1001000: c <= 9'b111000111;
				8'b111000: c <= 9'b110011110;
				8'b110001: c <= 9'b11001101;
				8'b1010111: c <= 9'b11;
				8'b1001110: c <= 9'b100000001;
				8'b1101010: c <= 9'b101000111;
				8'b1001001: c <= 9'b101001000;
				8'b1100000: c <= 9'b10110101;
				8'b110111: c <= 9'b11001101;
				8'b1011101: c <= 9'b1000000;
				8'b1011011: c <= 9'b10001111;
				8'b111001: c <= 9'b11101100;
				8'b1001010: c <= 9'b10101;
				8'b110011: c <= 9'b100110;
				8'b1101100: c <= 9'b1100100;
				8'b1110111: c <= 9'b110010011;
				8'b101011: c <= 9'b1001000;
				8'b1101011: c <= 9'b10001100;
				8'b111100: c <= 9'b10110010;
				8'b1000111: c <= 9'b110011001;
				8'b1011111: c <= 9'b100000010;
				8'b1110100: c <= 9'b11001;
				8'b101101: c <= 9'b100101010;
				8'b1010011: c <= 9'b1100110;
				8'b1100001: c <= 9'b100100;
				8'b110101: c <= 9'b10111000;
				8'b1000100: c <= 9'b10011010;
				8'b1010001: c <= 9'b101101011;
				8'b1010100: c <= 9'b110111110;
				8'b1100110: c <= 9'b100011000;
				8'b101010: c <= 9'b111101100;
				8'b1011110: c <= 9'b1101110;
				8'b1100111: c <= 9'b11100000;
				8'b1011010: c <= 9'b10110101;
				8'b1000010: c <= 9'b111101111;
				8'b111101: c <= 9'b110101001;
				8'b110000: c <= 9'b110110110;
				8'b111110: c <= 9'b11101100;
				8'b1100010: c <= 9'b1111000;
				8'b1110000: c <= 9'b10000111;
				8'b1101001: c <= 9'b1101;
				8'b1110011: c <= 9'b110101100;
				8'b1001100: c <= 9'b110100110;
				8'b100001: c <= 9'b110000000;
				8'b1000110: c <= 9'b100111001;
				8'b1110010: c <= 9'b100111100;
				8'b1010000: c <= 9'b111000011;
				8'b1111010: c <= 9'b101010110;
				8'b1010101: c <= 9'b110;
				8'b111011: c <= 9'b110000111;
				8'b1001101: c <= 9'b10110010;
				8'b111111: c <= 9'b100011100;
				8'b1101110: c <= 9'b10011111;
				8'b1111011: c <= 9'b11101;
				8'b1001011: c <= 9'b101110101;
				8'b1101111: c <= 9'b11110000;
				8'b1101000: c <= 9'b100010100;
				8'b101100: c <= 9'b10100;
				8'b100100: c <= 9'b100111010;
				8'b1111000: c <= 9'b101100100;
				8'b1000101: c <= 9'b1110001;
				8'b1011001: c <= 9'b111001111;
				8'b110100: c <= 9'b1111010;
				8'b1111001: c <= 9'b101111111;
				8'b1110001: c <= 9'b10110010;
				8'b1001111: c <= 9'b10100111;
				8'b1100101: c <= 9'b10101101;
				8'b1111110: c <= 9'b110110111;
				8'b1111100: c <= 9'b11100001;
				8'b1010110: c <= 9'b110010110;
				8'b110010: c <= 9'b100010111;
				8'b1101101: c <= 9'b1011001;
				8'b100011: c <= 9'b100111101;
				8'b1110101: c <= 9'b11;
				8'b1111101: c <= 9'b111100011;
				8'b101001: c <= 9'b110000011;
				8'b1010010: c <= 9'b111101000;
				8'b1011000: c <= 9'b101000011;
				8'b101110: c <= 9'b11100111;
				8'b1000001: c <= 9'b101110001;
				default: c <= 9'b0;
			endcase
			9'b10100101 : case(di)
				8'b1000011: c <= 9'b1;
				8'b101000: c <= 9'b1001011;
				8'b111010: c <= 9'b101001111;
				8'b110110: c <= 9'b1100011;
				8'b1100100: c <= 9'b100;
				8'b1000000: c <= 9'b111111110;
				8'b1110110: c <= 9'b100110111;
				8'b100101: c <= 9'b110010111;
				8'b101111: c <= 9'b101010;
				8'b100110: c <= 9'b11111101;
				8'b1100011: c <= 9'b1101111;
				8'b1001000: c <= 9'b110111110;
				8'b111000: c <= 9'b110011100;
				8'b110001: c <= 9'b110110111;
				8'b1010111: c <= 9'b11001100;
				8'b1001110: c <= 9'b11110011;
				8'b1101010: c <= 9'b10101101;
				8'b1001001: c <= 9'b111011110;
				8'b1100000: c <= 9'b10;
				8'b110111: c <= 9'b101001110;
				8'b1011101: c <= 9'b100000111;
				8'b1011011: c <= 9'b111111110;
				8'b111001: c <= 9'b110110000;
				8'b1001010: c <= 9'b101101111;
				8'b110011: c <= 9'b100011000;
				8'b1101100: c <= 9'b110110100;
				8'b1110111: c <= 9'b100001010;
				8'b101011: c <= 9'b100011001;
				8'b1101011: c <= 9'b11110100;
				8'b111100: c <= 9'b101000111;
				8'b1000111: c <= 9'b101010000;
				8'b1011111: c <= 9'b101010;
				8'b1110100: c <= 9'b10101001;
				8'b101101: c <= 9'b100001101;
				8'b1010011: c <= 9'b11111101;
				8'b1100001: c <= 9'b11100000;
				8'b110101: c <= 9'b1010110;
				8'b1000100: c <= 9'b101110;
				8'b1010001: c <= 9'b11010101;
				8'b1010100: c <= 9'b1101001;
				8'b1100110: c <= 9'b10001000;
				8'b101010: c <= 9'b11100001;
				8'b1011110: c <= 9'b11101011;
				8'b1100111: c <= 9'b11110000;
				8'b1011010: c <= 9'b1100;
				8'b1000010: c <= 9'b10001100;
				8'b111101: c <= 9'b1101000;
				8'b110000: c <= 9'b10010111;
				8'b111110: c <= 9'b100100010;
				8'b1100010: c <= 9'b11000100;
				8'b1110000: c <= 9'b101101100;
				8'b1101001: c <= 9'b10111001;
				8'b1110011: c <= 9'b1000101;
				8'b1001100: c <= 9'b10100101;
				8'b100001: c <= 9'b100111011;
				8'b1000110: c <= 9'b1001010;
				8'b1110010: c <= 9'b100000000;
				8'b1010000: c <= 9'b11010111;
				8'b1111010: c <= 9'b100110000;
				8'b1010101: c <= 9'b1101000;
				8'b111011: c <= 9'b111010111;
				8'b1001101: c <= 9'b10010000;
				8'b111111: c <= 9'b100000111;
				8'b1101110: c <= 9'b10111101;
				8'b1111011: c <= 9'b101011101;
				8'b1001011: c <= 9'b1100011;
				8'b1101111: c <= 9'b101110110;
				8'b1101000: c <= 9'b1;
				8'b101100: c <= 9'b111001110;
				8'b100100: c <= 9'b10101101;
				8'b1111000: c <= 9'b110001011;
				8'b1000101: c <= 9'b111100100;
				8'b1011001: c <= 9'b110001101;
				8'b110100: c <= 9'b1011000;
				8'b1111001: c <= 9'b10000101;
				8'b1110001: c <= 9'b111001010;
				8'b1001111: c <= 9'b110100101;
				8'b1100101: c <= 9'b110100001;
				8'b1111110: c <= 9'b110000010;
				8'b1111100: c <= 9'b101101;
				8'b1010110: c <= 9'b111010;
				8'b110010: c <= 9'b1110000;
				8'b1101101: c <= 9'b111000010;
				8'b100011: c <= 9'b10000000;
				8'b1110101: c <= 9'b1110111;
				8'b1111101: c <= 9'b111000100;
				8'b101001: c <= 9'b111101;
				8'b1010010: c <= 9'b1000010;
				8'b1011000: c <= 9'b101000011;
				8'b101110: c <= 9'b10001000;
				8'b1000001: c <= 9'b1001010;
				default: c <= 9'b0;
			endcase
			9'b1101111 : case(di)
				8'b1000011: c <= 9'b101100011;
				8'b101000: c <= 9'b101110100;
				8'b111010: c <= 9'b111001111;
				8'b110110: c <= 9'b101010100;
				8'b1100100: c <= 9'b1111011;
				8'b1000000: c <= 9'b11010001;
				8'b1110110: c <= 9'b111101101;
				8'b100101: c <= 9'b101010000;
				8'b101111: c <= 9'b11110;
				8'b100110: c <= 9'b10;
				8'b1100011: c <= 9'b101011001;
				8'b1001000: c <= 9'b10010011;
				8'b111000: c <= 9'b11101000;
				8'b110001: c <= 9'b101011111;
				8'b1010111: c <= 9'b10111001;
				8'b1001110: c <= 9'b111011;
				8'b1101010: c <= 9'b10100;
				8'b1001001: c <= 9'b110010100;
				8'b1100000: c <= 9'b101000;
				8'b110111: c <= 9'b101010010;
				8'b1011101: c <= 9'b1101001;
				8'b1011011: c <= 9'b110000110;
				8'b111001: c <= 9'b11100000;
				8'b1001010: c <= 9'b100001101;
				8'b110011: c <= 9'b10101;
				8'b1101100: c <= 9'b100001001;
				8'b1110111: c <= 9'b100100110;
				8'b101011: c <= 9'b10001010;
				8'b1101011: c <= 9'b100101;
				8'b111100: c <= 9'b110100100;
				8'b1000111: c <= 9'b100101010;
				8'b1011111: c <= 9'b110001010;
				8'b1110100: c <= 9'b11111101;
				8'b101101: c <= 9'b11100010;
				8'b1010011: c <= 9'b11010101;
				8'b1100001: c <= 9'b110101;
				8'b110101: c <= 9'b11100101;
				8'b1000100: c <= 9'b101101010;
				8'b1010001: c <= 9'b100001101;
				8'b1010100: c <= 9'b110100011;
				8'b1100110: c <= 9'b110101101;
				8'b101010: c <= 9'b101011;
				8'b1011110: c <= 9'b101111000;
				8'b1100111: c <= 9'b101101010;
				8'b1011010: c <= 9'b110010101;
				8'b1000010: c <= 9'b110111010;
				8'b111101: c <= 9'b101111110;
				8'b110000: c <= 9'b11000010;
				8'b111110: c <= 9'b111000;
				8'b1100010: c <= 9'b100000011;
				8'b1110000: c <= 9'b10011101;
				8'b1101001: c <= 9'b100011;
				8'b1110011: c <= 9'b10110001;
				8'b1001100: c <= 9'b10010110;
				8'b100001: c <= 9'b10100101;
				8'b1000110: c <= 9'b111011100;
				8'b1110010: c <= 9'b11110000;
				8'b1010000: c <= 9'b100110111;
				8'b1111010: c <= 9'b1111000;
				8'b1010101: c <= 9'b10011001;
				8'b111011: c <= 9'b111101000;
				8'b1001101: c <= 9'b110011111;
				8'b111111: c <= 9'b110101101;
				8'b1101110: c <= 9'b11110000;
				8'b1111011: c <= 9'b111111;
				8'b1001011: c <= 9'b111110001;
				8'b1101111: c <= 9'b11010000;
				8'b1101000: c <= 9'b111101001;
				8'b101100: c <= 9'b110101111;
				8'b100100: c <= 9'b111011100;
				8'b1111000: c <= 9'b11110110;
				8'b1000101: c <= 9'b11001101;
				8'b1011001: c <= 9'b10000011;
				8'b110100: c <= 9'b1110101;
				8'b1111001: c <= 9'b101111001;
				8'b1110001: c <= 9'b10010000;
				8'b1001111: c <= 9'b1101100;
				8'b1100101: c <= 9'b111000;
				8'b1111110: c <= 9'b111101010;
				8'b1111100: c <= 9'b100000010;
				8'b1010110: c <= 9'b11100000;
				8'b110010: c <= 9'b110010100;
				8'b1101101: c <= 9'b100101000;
				8'b100011: c <= 9'b11001010;
				8'b1110101: c <= 9'b110100101;
				8'b1111101: c <= 9'b110111011;
				8'b101001: c <= 9'b100011000;
				8'b1010010: c <= 9'b110111001;
				8'b1011000: c <= 9'b101100111;
				8'b101110: c <= 9'b100111000;
				8'b1000001: c <= 9'b11001111;
				default: c <= 9'b0;
			endcase
			9'b10101001 : case(di)
				8'b1000011: c <= 9'b101010011;
				8'b101000: c <= 9'b10111010;
				8'b111010: c <= 9'b111000100;
				8'b110110: c <= 9'b101100011;
				8'b1100100: c <= 9'b11001001;
				8'b1000000: c <= 9'b111010000;
				8'b1110110: c <= 9'b100100111;
				8'b100101: c <= 9'b101011000;
				8'b101111: c <= 9'b10010110;
				8'b100110: c <= 9'b110110011;
				8'b1100011: c <= 9'b10011;
				8'b1001000: c <= 9'b100011101;
				8'b111000: c <= 9'b100000101;
				8'b110001: c <= 9'b101101010;
				8'b1010111: c <= 9'b1011011;
				8'b1001110: c <= 9'b1001;
				8'b1101010: c <= 9'b11000110;
				8'b1001001: c <= 9'b100011000;
				8'b1100000: c <= 9'b101100001;
				8'b110111: c <= 9'b1011011;
				8'b1011101: c <= 9'b1001110;
				8'b1011011: c <= 9'b111010111;
				8'b111001: c <= 9'b10010011;
				8'b1001010: c <= 9'b1111001;
				8'b110011: c <= 9'b1100;
				8'b1101100: c <= 9'b111110001;
				8'b1110111: c <= 9'b101110000;
				8'b101011: c <= 9'b1110100;
				8'b1101011: c <= 9'b100111;
				8'b111100: c <= 9'b1101111;
				8'b1000111: c <= 9'b100101111;
				8'b1011111: c <= 9'b100001101;
				8'b1110100: c <= 9'b10110100;
				8'b101101: c <= 9'b1111;
				8'b1010011: c <= 9'b100000011;
				8'b1100001: c <= 9'b100110100;
				8'b110101: c <= 9'b10010111;
				8'b1000100: c <= 9'b10010011;
				8'b1010001: c <= 9'b1000110;
				8'b1010100: c <= 9'b101100;
				8'b1100110: c <= 9'b101100111;
				8'b101010: c <= 9'b10010;
				8'b1011110: c <= 9'b100101111;
				8'b1100111: c <= 9'b10100111;
				8'b1011010: c <= 9'b100011001;
				8'b1000010: c <= 9'b101000011;
				8'b111101: c <= 9'b100011;
				8'b110000: c <= 9'b110001000;
				8'b111110: c <= 9'b10100;
				8'b1100010: c <= 9'b100010;
				8'b1110000: c <= 9'b111101110;
				8'b1101001: c <= 9'b110000110;
				8'b1110011: c <= 9'b100010111;
				8'b1001100: c <= 9'b100001011;
				8'b100001: c <= 9'b111111011;
				8'b1000110: c <= 9'b10000000;
				8'b1110010: c <= 9'b110111;
				8'b1010000: c <= 9'b11101111;
				8'b1111010: c <= 9'b111000110;
				8'b1010101: c <= 9'b100100101;
				8'b111011: c <= 9'b1010010;
				8'b1001101: c <= 9'b110010101;
				8'b111111: c <= 9'b10100011;
				8'b1101110: c <= 9'b10101111;
				8'b1111011: c <= 9'b1011110;
				8'b1001011: c <= 9'b10010111;
				8'b1101111: c <= 9'b101101000;
				8'b1101000: c <= 9'b100011100;
				8'b101100: c <= 9'b1001001;
				8'b100100: c <= 9'b1110011;
				8'b1111000: c <= 9'b101110;
				8'b1000101: c <= 9'b10001001;
				8'b1011001: c <= 9'b110111000;
				8'b110100: c <= 9'b110001;
				8'b1111001: c <= 9'b1101100;
				8'b1110001: c <= 9'b1001100;
				8'b1001111: c <= 9'b1101111;
				8'b1100101: c <= 9'b111101010;
				8'b1111110: c <= 9'b101011;
				8'b1111100: c <= 9'b100100001;
				8'b1010110: c <= 9'b111;
				8'b110010: c <= 9'b111100101;
				8'b1101101: c <= 9'b110111001;
				8'b100011: c <= 9'b100111010;
				8'b1110101: c <= 9'b1011000;
				8'b1111101: c <= 9'b111100110;
				8'b101001: c <= 9'b111101111;
				8'b1010010: c <= 9'b1001101;
				8'b1011000: c <= 9'b11010010;
				8'b101110: c <= 9'b110101001;
				8'b1000001: c <= 9'b11011101;
				default: c <= 9'b0;
			endcase
			9'b101011001 : case(di)
				8'b1000011: c <= 9'b11011000;
				8'b101000: c <= 9'b1011000;
				8'b111010: c <= 9'b11000110;
				8'b110110: c <= 9'b11000001;
				8'b1100100: c <= 9'b101011010;
				8'b1000000: c <= 9'b11000111;
				8'b1110110: c <= 9'b110001;
				8'b100101: c <= 9'b1100010;
				8'b101111: c <= 9'b110011;
				8'b100110: c <= 9'b111000111;
				8'b1100011: c <= 9'b111100000;
				8'b1001000: c <= 9'b101101011;
				8'b111000: c <= 9'b10110010;
				8'b110001: c <= 9'b111101111;
				8'b1010111: c <= 9'b111011;
				8'b1001110: c <= 9'b10010101;
				8'b1101010: c <= 9'b110100111;
				8'b1001001: c <= 9'b1001011;
				8'b1100000: c <= 9'b111000100;
				8'b110111: c <= 9'b10011100;
				8'b1011101: c <= 9'b100001010;
				8'b1011011: c <= 9'b11100010;
				8'b111001: c <= 9'b111110110;
				8'b1001010: c <= 9'b100010;
				8'b110011: c <= 9'b1101110;
				8'b1101100: c <= 9'b101011;
				8'b1110111: c <= 9'b1101010;
				8'b101011: c <= 9'b101010010;
				8'b1101011: c <= 9'b100100110;
				8'b111100: c <= 9'b111010110;
				8'b1000111: c <= 9'b101000111;
				8'b1011111: c <= 9'b10110;
				8'b1110100: c <= 9'b111101110;
				8'b101101: c <= 9'b10001100;
				8'b1010011: c <= 9'b111111110;
				8'b1100001: c <= 9'b111011;
				8'b110101: c <= 9'b10100101;
				8'b1000100: c <= 9'b1101101;
				8'b1010001: c <= 9'b111111000;
				8'b1010100: c <= 9'b11110000;
				8'b1100110: c <= 9'b101011011;
				8'b101010: c <= 9'b111010010;
				8'b1011110: c <= 9'b11100100;
				8'b1100111: c <= 9'b110101001;
				8'b1011010: c <= 9'b11110011;
				8'b1000010: c <= 9'b111000101;
				8'b111101: c <= 9'b11101000;
				8'b110000: c <= 9'b1101100;
				8'b111110: c <= 9'b1110001;
				8'b1100010: c <= 9'b10011010;
				8'b1110000: c <= 9'b100100011;
				8'b1101001: c <= 9'b10101111;
				8'b1110011: c <= 9'b101100010;
				8'b1001100: c <= 9'b110011010;
				8'b100001: c <= 9'b101010001;
				8'b1000110: c <= 9'b11101000;
				8'b1110010: c <= 9'b100111010;
				8'b1010000: c <= 9'b110011101;
				8'b1111010: c <= 9'b101111000;
				8'b1010101: c <= 9'b111001110;
				8'b111011: c <= 9'b100011000;
				8'b1001101: c <= 9'b100001;
				8'b111111: c <= 9'b110011100;
				8'b1101110: c <= 9'b10110110;
				8'b1111011: c <= 9'b100010100;
				8'b1001011: c <= 9'b1001110;
				8'b1101111: c <= 9'b110100;
				8'b1101000: c <= 9'b101000010;
				8'b101100: c <= 9'b11011010;
				8'b100100: c <= 9'b110000011;
				8'b1111000: c <= 9'b11100;
				8'b1000101: c <= 9'b11100010;
				8'b1011001: c <= 9'b11110100;
				8'b110100: c <= 9'b1111101;
				8'b1111001: c <= 9'b1011100;
				8'b1110001: c <= 9'b101011111;
				8'b1001111: c <= 9'b110101001;
				8'b1100101: c <= 9'b111011001;
				8'b1111110: c <= 9'b111101;
				8'b1111100: c <= 9'b10111110;
				8'b1010110: c <= 9'b1110101;
				8'b110010: c <= 9'b11110011;
				8'b1101101: c <= 9'b11101000;
				8'b100011: c <= 9'b111000110;
				8'b1110101: c <= 9'b110010101;
				8'b1111101: c <= 9'b110000101;
				8'b101001: c <= 9'b101110110;
				8'b1010010: c <= 9'b100110000;
				8'b1011000: c <= 9'b111010010;
				8'b101110: c <= 9'b11111010;
				8'b1000001: c <= 9'b110101100;
				default: c <= 9'b0;
			endcase
			9'b11010000 : case(di)
				8'b1000011: c <= 9'b111100;
				8'b101000: c <= 9'b101110110;
				8'b111010: c <= 9'b110110101;
				8'b110110: c <= 9'b10001101;
				8'b1100100: c <= 9'b1101100;
				8'b1000000: c <= 9'b111010000;
				8'b1110110: c <= 9'b11010010;
				8'b100101: c <= 9'b10100010;
				8'b101111: c <= 9'b110101;
				8'b100110: c <= 9'b101010000;
				8'b1100011: c <= 9'b110101011;
				8'b1001000: c <= 9'b101100101;
				8'b111000: c <= 9'b110101110;
				8'b110001: c <= 9'b101000110;
				8'b1010111: c <= 9'b11000001;
				8'b1001110: c <= 9'b110001001;
				8'b1101010: c <= 9'b101111001;
				8'b1001001: c <= 9'b111011011;
				8'b1100000: c <= 9'b110010101;
				8'b110111: c <= 9'b101111110;
				8'b1011101: c <= 9'b1111110;
				8'b1011011: c <= 9'b110000011;
				8'b111001: c <= 9'b10011000;
				8'b1001010: c <= 9'b101;
				8'b110011: c <= 9'b10;
				8'b1101100: c <= 9'b10000011;
				8'b1110111: c <= 9'b110000001;
				8'b101011: c <= 9'b11100011;
				8'b1101011: c <= 9'b11010001;
				8'b111100: c <= 9'b110011100;
				8'b1000111: c <= 9'b1101000;
				8'b1011111: c <= 9'b100010100;
				8'b1110100: c <= 9'b111111000;
				8'b101101: c <= 9'b101101111;
				8'b1010011: c <= 9'b11111100;
				8'b1100001: c <= 9'b11001101;
				8'b110101: c <= 9'b1010110;
				8'b1000100: c <= 9'b11011001;
				8'b1010001: c <= 9'b110110101;
				8'b1010100: c <= 9'b1010111;
				8'b1100110: c <= 9'b100101101;
				8'b101010: c <= 9'b10001110;
				8'b1011110: c <= 9'b110000110;
				8'b1100111: c <= 9'b1000100;
				8'b1011010: c <= 9'b1100111;
				8'b1000010: c <= 9'b101100011;
				8'b111101: c <= 9'b111011;
				8'b110000: c <= 9'b10010;
				8'b111110: c <= 9'b110101010;
				8'b1100010: c <= 9'b10010000;
				8'b1110000: c <= 9'b1111;
				8'b1101001: c <= 9'b10000010;
				8'b1110011: c <= 9'b111101101;
				8'b1001100: c <= 9'b10101100;
				8'b100001: c <= 9'b100001101;
				8'b1000110: c <= 9'b1000001;
				8'b1110010: c <= 9'b111000011;
				8'b1010000: c <= 9'b110101;
				8'b1111010: c <= 9'b111011110;
				8'b1010101: c <= 9'b110011101;
				8'b111011: c <= 9'b100100001;
				8'b1001101: c <= 9'b1110100;
				8'b111111: c <= 9'b11110001;
				8'b1101110: c <= 9'b101010100;
				8'b1111011: c <= 9'b100110;
				8'b1001011: c <= 9'b100100011;
				8'b1101111: c <= 9'b101101010;
				8'b1101000: c <= 9'b110100110;
				8'b101100: c <= 9'b11001100;
				8'b100100: c <= 9'b100001001;
				8'b1111000: c <= 9'b110101100;
				8'b1000101: c <= 9'b101011011;
				8'b1011001: c <= 9'b1001000;
				8'b110100: c <= 9'b110100101;
				8'b1111001: c <= 9'b101100;
				8'b1110001: c <= 9'b101111010;
				8'b1001111: c <= 9'b110010010;
				8'b1100101: c <= 9'b101100100;
				8'b1111110: c <= 9'b110011100;
				8'b1111100: c <= 9'b100110100;
				8'b1010110: c <= 9'b110100001;
				8'b110010: c <= 9'b111110000;
				8'b1101101: c <= 9'b11100110;
				8'b100011: c <= 9'b10101101;
				8'b1110101: c <= 9'b110101101;
				8'b1111101: c <= 9'b11110011;
				8'b101001: c <= 9'b110110;
				8'b1010010: c <= 9'b101001011;
				8'b1011000: c <= 9'b1000100;
				8'b101110: c <= 9'b10010001;
				8'b1000001: c <= 9'b1110;
				default: c <= 9'b0;
			endcase
			9'b1010111 : case(di)
				8'b1000011: c <= 9'b10110001;
				8'b101000: c <= 9'b111110000;
				8'b111010: c <= 9'b111111101;
				8'b110110: c <= 9'b111001010;
				8'b1100100: c <= 9'b10010100;
				8'b1000000: c <= 9'b111001111;
				8'b1110110: c <= 9'b11001111;
				8'b100101: c <= 9'b101;
				8'b101111: c <= 9'b1010010;
				8'b100110: c <= 9'b110000001;
				8'b1100011: c <= 9'b101001111;
				8'b1001000: c <= 9'b10111100;
				8'b111000: c <= 9'b100110010;
				8'b110001: c <= 9'b110010;
				8'b1010111: c <= 9'b111101100;
				8'b1001110: c <= 9'b1000110;
				8'b1101010: c <= 9'b110111;
				8'b1001001: c <= 9'b1011100;
				8'b1100000: c <= 9'b1111010;
				8'b110111: c <= 9'b11111010;
				8'b1011101: c <= 9'b1111101;
				8'b1011011: c <= 9'b100101001;
				8'b111001: c <= 9'b110101111;
				8'b1001010: c <= 9'b100100000;
				8'b110011: c <= 9'b11111110;
				8'b1101100: c <= 9'b100010000;
				8'b1110111: c <= 9'b101101101;
				8'b101011: c <= 9'b10111101;
				8'b1101011: c <= 9'b11101000;
				8'b111100: c <= 9'b11000010;
				8'b1000111: c <= 9'b11110011;
				8'b1011111: c <= 9'b100010;
				8'b1110100: c <= 9'b111010100;
				8'b101101: c <= 9'b100011111;
				8'b1010011: c <= 9'b100000101;
				8'b1100001: c <= 9'b10100101;
				8'b110101: c <= 9'b101110101;
				8'b1000100: c <= 9'b1001011;
				8'b1010001: c <= 9'b111011011;
				8'b1010100: c <= 9'b1101001;
				8'b1100110: c <= 9'b110011000;
				8'b101010: c <= 9'b100001;
				8'b1011110: c <= 9'b11011;
				8'b1100111: c <= 9'b100000110;
				8'b1011010: c <= 9'b100000011;
				8'b1000010: c <= 9'b110001011;
				8'b111101: c <= 9'b101111001;
				8'b110000: c <= 9'b11010101;
				8'b111110: c <= 9'b111111000;
				8'b1100010: c <= 9'b110110000;
				8'b1110000: c <= 9'b1101;
				8'b1101001: c <= 9'b111101;
				8'b1110011: c <= 9'b100001101;
				8'b1001100: c <= 9'b111110001;
				8'b100001: c <= 9'b11111001;
				8'b1000110: c <= 9'b110;
				8'b1110010: c <= 9'b111010111;
				8'b1010000: c <= 9'b101110101;
				8'b1111010: c <= 9'b110101101;
				8'b1010101: c <= 9'b100110111;
				8'b111011: c <= 9'b1001110;
				8'b1001101: c <= 9'b110100010;
				8'b111111: c <= 9'b11100;
				8'b1101110: c <= 9'b100110010;
				8'b1111011: c <= 9'b110011110;
				8'b1001011: c <= 9'b101000010;
				8'b1101111: c <= 9'b110001101;
				8'b1101000: c <= 9'b110001000;
				8'b101100: c <= 9'b111100010;
				8'b100100: c <= 9'b100101110;
				8'b1111000: c <= 9'b11001100;
				8'b1000101: c <= 9'b101101110;
				8'b1011001: c <= 9'b111100010;
				8'b110100: c <= 9'b110000111;
				8'b1111001: c <= 9'b100110111;
				8'b1110001: c <= 9'b10101110;
				8'b1001111: c <= 9'b110100;
				8'b1100101: c <= 9'b1100101;
				8'b1111110: c <= 9'b110110101;
				8'b1111100: c <= 9'b110001101;
				8'b1010110: c <= 9'b1100001;
				8'b110010: c <= 9'b110101;
				8'b1101101: c <= 9'b111110000;
				8'b100011: c <= 9'b11000011;
				8'b1110101: c <= 9'b100110110;
				8'b1111101: c <= 9'b11011110;
				8'b101001: c <= 9'b110011001;
				8'b1010010: c <= 9'b11010001;
				8'b1011000: c <= 9'b111010000;
				8'b101110: c <= 9'b1111;
				8'b1000001: c <= 9'b101011;
				default: c <= 9'b0;
			endcase
			9'b111111 : case(di)
				8'b1000011: c <= 9'b11110100;
				8'b101000: c <= 9'b1010000;
				8'b111010: c <= 9'b100001;
				8'b110110: c <= 9'b101100010;
				8'b1100100: c <= 9'b100101010;
				8'b1000000: c <= 9'b11000;
				8'b1110110: c <= 9'b11010001;
				8'b100101: c <= 9'b101010101;
				8'b101111: c <= 9'b10101111;
				8'b100110: c <= 9'b1100100;
				8'b1100011: c <= 9'b110000010;
				8'b1001000: c <= 9'b100100010;
				8'b111000: c <= 9'b111111011;
				8'b110001: c <= 9'b11110;
				8'b1010111: c <= 9'b11110;
				8'b1001110: c <= 9'b10010100;
				8'b1101010: c <= 9'b1111100;
				8'b1001001: c <= 9'b1011001;
				8'b1100000: c <= 9'b111110101;
				8'b110111: c <= 9'b110011000;
				8'b1011101: c <= 9'b11011110;
				8'b1011011: c <= 9'b11100110;
				8'b111001: c <= 9'b11011110;
				8'b1001010: c <= 9'b10111000;
				8'b110011: c <= 9'b10011000;
				8'b1101100: c <= 9'b100001001;
				8'b1110111: c <= 9'b111000010;
				8'b101011: c <= 9'b100101;
				8'b1101011: c <= 9'b11101100;
				8'b111100: c <= 9'b101010010;
				8'b1000111: c <= 9'b1011011;
				8'b1011111: c <= 9'b101011001;
				8'b1110100: c <= 9'b10110110;
				8'b101101: c <= 9'b100111011;
				8'b1010011: c <= 9'b1001110;
				8'b1100001: c <= 9'b100001100;
				8'b110101: c <= 9'b11001111;
				8'b1000100: c <= 9'b1100011;
				8'b1010001: c <= 9'b10011100;
				8'b1010100: c <= 9'b11111000;
				8'b1100110: c <= 9'b1100101;
				8'b101010: c <= 9'b100001;
				8'b1011110: c <= 9'b1111010;
				8'b1100111: c <= 9'b1000010;
				8'b1011010: c <= 9'b110111110;
				8'b1000010: c <= 9'b11111011;
				8'b111101: c <= 9'b10101101;
				8'b110000: c <= 9'b100011111;
				8'b111110: c <= 9'b101000001;
				8'b1100010: c <= 9'b100001001;
				8'b1110000: c <= 9'b1100101;
				8'b1101001: c <= 9'b111001;
				8'b1110011: c <= 9'b11001110;
				8'b1001100: c <= 9'b101010010;
				8'b100001: c <= 9'b101110101;
				8'b1000110: c <= 9'b111001000;
				8'b1110010: c <= 9'b100101011;
				8'b1010000: c <= 9'b1100001;
				8'b1111010: c <= 9'b100011001;
				8'b1010101: c <= 9'b110110101;
				8'b111011: c <= 9'b110101010;
				8'b1001101: c <= 9'b110110110;
				8'b111111: c <= 9'b11110111;
				8'b1101110: c <= 9'b111101100;
				8'b1111011: c <= 9'b111001110;
				8'b1001011: c <= 9'b1001110;
				8'b1101111: c <= 9'b100010000;
				8'b1101000: c <= 9'b100;
				8'b101100: c <= 9'b11011000;
				8'b100100: c <= 9'b10100011;
				8'b1111000: c <= 9'b1110011;
				8'b1000101: c <= 9'b110000001;
				8'b1011001: c <= 9'b11010000;
				8'b110100: c <= 9'b1110111;
				8'b1111001: c <= 9'b111011011;
				8'b1110001: c <= 9'b100100010;
				8'b1001111: c <= 9'b101010101;
				8'b1100101: c <= 9'b111101110;
				8'b1111110: c <= 9'b101;
				8'b1111100: c <= 9'b110110010;
				8'b1010110: c <= 9'b101110000;
				8'b110010: c <= 9'b10100000;
				8'b1101101: c <= 9'b10000000;
				8'b100011: c <= 9'b10001110;
				8'b1110101: c <= 9'b11100010;
				8'b1111101: c <= 9'b100010001;
				8'b101001: c <= 9'b101011111;
				8'b1010010: c <= 9'b111001;
				8'b1011000: c <= 9'b10101001;
				8'b101110: c <= 9'b10101011;
				8'b1000001: c <= 9'b11000011;
				default: c <= 9'b0;
			endcase
			9'b10000010 : case(di)
				8'b1000011: c <= 9'b1101111;
				8'b101000: c <= 9'b101010010;
				8'b111010: c <= 9'b110001110;
				8'b110110: c <= 9'b100010001;
				8'b1100100: c <= 9'b111011110;
				8'b1000000: c <= 9'b111100011;
				8'b1110110: c <= 9'b110110000;
				8'b100101: c <= 9'b11010;
				8'b101111: c <= 9'b111111101;
				8'b100110: c <= 9'b1011110;
				8'b1100011: c <= 9'b11111010;
				8'b1001000: c <= 9'b1010000;
				8'b111000: c <= 9'b110011111;
				8'b110001: c <= 9'b101010100;
				8'b1010111: c <= 9'b1000;
				8'b1001110: c <= 9'b110000110;
				8'b1101010: c <= 9'b1101010;
				8'b1001001: c <= 9'b1001011;
				8'b1100000: c <= 9'b101100001;
				8'b110111: c <= 9'b100100110;
				8'b1011101: c <= 9'b100101111;
				8'b1011011: c <= 9'b110011100;
				8'b111001: c <= 9'b10101000;
				8'b1001010: c <= 9'b100010000;
				8'b110011: c <= 9'b110110110;
				8'b1101100: c <= 9'b101111010;
				8'b1110111: c <= 9'b11111011;
				8'b101011: c <= 9'b100001101;
				8'b1101011: c <= 9'b11110111;
				8'b111100: c <= 9'b101111010;
				8'b1000111: c <= 9'b110001101;
				8'b1011111: c <= 9'b101101011;
				8'b1110100: c <= 9'b101010010;
				8'b101101: c <= 9'b1100001;
				8'b1010011: c <= 9'b111100110;
				8'b1100001: c <= 9'b100101010;
				8'b110101: c <= 9'b111010010;
				8'b1000100: c <= 9'b111110000;
				8'b1010001: c <= 9'b110011101;
				8'b1010100: c <= 9'b100111010;
				8'b1100110: c <= 9'b11110000;
				8'b101010: c <= 9'b101100100;
				8'b1011110: c <= 9'b101010100;
				8'b1100111: c <= 9'b101010101;
				8'b1011010: c <= 9'b10110010;
				8'b1000010: c <= 9'b1101000;
				8'b111101: c <= 9'b100101110;
				8'b110000: c <= 9'b1001;
				8'b111110: c <= 9'b110101011;
				8'b1100010: c <= 9'b11110110;
				8'b1110000: c <= 9'b101111000;
				8'b1101001: c <= 9'b1001;
				8'b1110011: c <= 9'b11101111;
				8'b1001100: c <= 9'b101001111;
				8'b100001: c <= 9'b111111000;
				8'b1000110: c <= 9'b100100001;
				8'b1110010: c <= 9'b101010000;
				8'b1010000: c <= 9'b111011011;
				8'b1111010: c <= 9'b110010101;
				8'b1010101: c <= 9'b100000000;
				8'b111011: c <= 9'b101110010;
				8'b1001101: c <= 9'b1010011;
				8'b111111: c <= 9'b11100011;
				8'b1101110: c <= 9'b101011010;
				8'b1111011: c <= 9'b110111111;
				8'b1001011: c <= 9'b110100;
				8'b1101111: c <= 9'b100111;
				8'b1101000: c <= 9'b10000000;
				8'b101100: c <= 9'b110110010;
				8'b100100: c <= 9'b110111111;
				8'b1111000: c <= 9'b111101010;
				8'b1000101: c <= 9'b10010100;
				8'b1011001: c <= 9'b1000010;
				8'b110100: c <= 9'b11100100;
				8'b1111001: c <= 9'b100010111;
				8'b1110001: c <= 9'b111101111;
				8'b1001111: c <= 9'b10011101;
				8'b1100101: c <= 9'b10100010;
				8'b1111110: c <= 9'b101111010;
				8'b1111100: c <= 9'b111111101;
				8'b1010110: c <= 9'b111101;
				8'b110010: c <= 9'b100110011;
				8'b1101101: c <= 9'b10000110;
				8'b100011: c <= 9'b111000010;
				8'b1110101: c <= 9'b10000110;
				8'b1111101: c <= 9'b101011011;
				8'b101001: c <= 9'b100;
				8'b1010010: c <= 9'b110100111;
				8'b1011000: c <= 9'b1010111;
				8'b101110: c <= 9'b10011001;
				8'b1000001: c <= 9'b1111000;
				default: c <= 9'b0;
			endcase
			9'b111111001 : case(di)
				8'b1000011: c <= 9'b111001000;
				8'b101000: c <= 9'b111010;
				8'b111010: c <= 9'b100010111;
				8'b110110: c <= 9'b101010111;
				8'b1100100: c <= 9'b10001100;
				8'b1000000: c <= 9'b110000111;
				8'b1110110: c <= 9'b1100001;
				8'b100101: c <= 9'b100001011;
				8'b101111: c <= 9'b100010;
				8'b100110: c <= 9'b11001111;
				8'b1100011: c <= 9'b111101;
				8'b1001000: c <= 9'b1011111;
				8'b111000: c <= 9'b111011001;
				8'b110001: c <= 9'b110010010;
				8'b1010111: c <= 9'b100111111;
				8'b1001110: c <= 9'b111000011;
				8'b1101010: c <= 9'b101100111;
				8'b1001001: c <= 9'b11100;
				8'b1100000: c <= 9'b110110110;
				8'b110111: c <= 9'b10101011;
				8'b1011101: c <= 9'b10111111;
				8'b1011011: c <= 9'b11101000;
				8'b111001: c <= 9'b1001100;
				8'b1001010: c <= 9'b1101001;
				8'b110011: c <= 9'b1000001;
				8'b1101100: c <= 9'b101100011;
				8'b1110111: c <= 9'b1101001;
				8'b101011: c <= 9'b101101000;
				8'b1101011: c <= 9'b101011011;
				8'b111100: c <= 9'b101011110;
				8'b1000111: c <= 9'b101011111;
				8'b1011111: c <= 9'b110011;
				8'b1110100: c <= 9'b101110111;
				8'b101101: c <= 9'b101100000;
				8'b1010011: c <= 9'b11011101;
				8'b1100001: c <= 9'b10000101;
				8'b110101: c <= 9'b111110101;
				8'b1000100: c <= 9'b101110111;
				8'b1010001: c <= 9'b110000;
				8'b1010100: c <= 9'b1101100;
				8'b1100110: c <= 9'b11110101;
				8'b101010: c <= 9'b11100100;
				8'b1011110: c <= 9'b1101000;
				8'b1100111: c <= 9'b1100100;
				8'b1011010: c <= 9'b1111;
				8'b1000010: c <= 9'b110101101;
				8'b111101: c <= 9'b11000110;
				8'b110000: c <= 9'b11110001;
				8'b111110: c <= 9'b110011111;
				8'b1100010: c <= 9'b1011001;
				8'b1110000: c <= 9'b111100011;
				8'b1101001: c <= 9'b10110010;
				8'b1110011: c <= 9'b100001011;
				8'b1001100: c <= 9'b101100010;
				8'b100001: c <= 9'b10110010;
				8'b1000110: c <= 9'b1010000;
				8'b1110010: c <= 9'b110000111;
				8'b1010000: c <= 9'b110100101;
				8'b1111010: c <= 9'b110011100;
				8'b1010101: c <= 9'b110001010;
				8'b111011: c <= 9'b11101001;
				8'b1001101: c <= 9'b1111001;
				8'b111111: c <= 9'b101110101;
				8'b1101110: c <= 9'b110101110;
				8'b1111011: c <= 9'b101010;
				8'b1001011: c <= 9'b100011;
				8'b1101111: c <= 9'b100000010;
				8'b1101000: c <= 9'b110011101;
				8'b101100: c <= 9'b10001110;
				8'b100100: c <= 9'b111000010;
				8'b1111000: c <= 9'b11010;
				8'b1000101: c <= 9'b1100001;
				8'b1011001: c <= 9'b101;
				8'b110100: c <= 9'b100101011;
				8'b1111001: c <= 9'b101010111;
				8'b1110001: c <= 9'b110111111;
				8'b1001111: c <= 9'b11110;
				8'b1100101: c <= 9'b100101;
				8'b1111110: c <= 9'b101001110;
				8'b1111100: c <= 9'b101110;
				8'b1010110: c <= 9'b100111101;
				8'b110010: c <= 9'b10100;
				8'b1101101: c <= 9'b10110011;
				8'b100011: c <= 9'b101010110;
				8'b1110101: c <= 9'b101011;
				8'b1111101: c <= 9'b10101100;
				8'b101001: c <= 9'b111001101;
				8'b1010010: c <= 9'b100011111;
				8'b1011000: c <= 9'b10001110;
				8'b101110: c <= 9'b1110100;
				8'b1000001: c <= 9'b10100110;
				default: c <= 9'b0;
			endcase
			9'b100100111 : case(di)
				8'b1000011: c <= 9'b10100;
				8'b101000: c <= 9'b10000010;
				8'b111010: c <= 9'b110011110;
				8'b110110: c <= 9'b1110100;
				8'b1100100: c <= 9'b101100010;
				8'b1000000: c <= 9'b111111111;
				8'b1110110: c <= 9'b100100101;
				8'b100101: c <= 9'b10001011;
				8'b101111: c <= 9'b1101;
				8'b100110: c <= 9'b11010010;
				8'b1100011: c <= 9'b100100101;
				8'b1001000: c <= 9'b111010;
				8'b111000: c <= 9'b111001111;
				8'b110001: c <= 9'b1110111;
				8'b1010111: c <= 9'b1101100;
				8'b1001110: c <= 9'b11001111;
				8'b1101010: c <= 9'b101010011;
				8'b1001001: c <= 9'b101110011;
				8'b1100000: c <= 9'b110100010;
				8'b110111: c <= 9'b111001100;
				8'b1011101: c <= 9'b111011111;
				8'b1011011: c <= 9'b100010111;
				8'b111001: c <= 9'b110001001;
				8'b1001010: c <= 9'b1100100;
				8'b110011: c <= 9'b1010110;
				8'b1101100: c <= 9'b101010;
				8'b1110111: c <= 9'b101110000;
				8'b101011: c <= 9'b101001000;
				8'b1101011: c <= 9'b10011101;
				8'b111100: c <= 9'b1110;
				8'b1000111: c <= 9'b111111;
				8'b1011111: c <= 9'b101010000;
				8'b1110100: c <= 9'b11000110;
				8'b101101: c <= 9'b110101101;
				8'b1010011: c <= 9'b1010000;
				8'b1100001: c <= 9'b10000000;
				8'b110101: c <= 9'b101110101;
				8'b1000100: c <= 9'b10111010;
				8'b1010001: c <= 9'b11011010;
				8'b1010100: c <= 9'b100010;
				8'b1100110: c <= 9'b110010101;
				8'b101010: c <= 9'b110011100;
				8'b1011110: c <= 9'b110101111;
				8'b1100111: c <= 9'b111111110;
				8'b1011010: c <= 9'b10010111;
				8'b1000010: c <= 9'b101000101;
				8'b111101: c <= 9'b110110110;
				8'b110000: c <= 9'b10010110;
				8'b111110: c <= 9'b111101111;
				8'b1100010: c <= 9'b10101011;
				8'b1110000: c <= 9'b11101100;
				8'b1101001: c <= 9'b1111;
				8'b1110011: c <= 9'b111000011;
				8'b1001100: c <= 9'b111001000;
				8'b100001: c <= 9'b100001111;
				8'b1000110: c <= 9'b11110;
				8'b1110010: c <= 9'b1011110;
				8'b1010000: c <= 9'b101000011;
				8'b1111010: c <= 9'b10001101;
				8'b1010101: c <= 9'b101110110;
				8'b111011: c <= 9'b11110000;
				8'b1001101: c <= 9'b100100000;
				8'b111111: c <= 9'b10001010;
				8'b1101110: c <= 9'b111001111;
				8'b1111011: c <= 9'b111000101;
				8'b1001011: c <= 9'b11011;
				8'b1101111: c <= 9'b10000111;
				8'b1101000: c <= 9'b10111111;
				8'b101100: c <= 9'b101011010;
				8'b100100: c <= 9'b110110110;
				8'b1111000: c <= 9'b110100100;
				8'b1000101: c <= 9'b1010111;
				8'b1011001: c <= 9'b10100011;
				8'b110100: c <= 9'b100101;
				8'b1111001: c <= 9'b111000000;
				8'b1110001: c <= 9'b10100111;
				8'b1001111: c <= 9'b100000010;
				8'b1100101: c <= 9'b1101010;
				8'b1111110: c <= 9'b100111010;
				8'b1111100: c <= 9'b100001111;
				8'b1010110: c <= 9'b10111010;
				8'b110010: c <= 9'b110010010;
				8'b1101101: c <= 9'b100100011;
				8'b100011: c <= 9'b1000101;
				8'b1110101: c <= 9'b10001111;
				8'b1111101: c <= 9'b100010110;
				8'b101001: c <= 9'b100010000;
				8'b1010010: c <= 9'b11101111;
				8'b1011000: c <= 9'b10001000;
				8'b101110: c <= 9'b101110001;
				8'b1000001: c <= 9'b101110101;
				default: c <= 9'b0;
			endcase
			9'b110101011 : case(di)
				8'b1000011: c <= 9'b100101010;
				8'b101000: c <= 9'b11110;
				8'b111010: c <= 9'b110001100;
				8'b110110: c <= 9'b100101001;
				8'b1100100: c <= 9'b111001;
				8'b1000000: c <= 9'b111000;
				8'b1110110: c <= 9'b11000010;
				8'b100101: c <= 9'b101100;
				8'b101111: c <= 9'b100001101;
				8'b100110: c <= 9'b1110001;
				8'b1100011: c <= 9'b110100111;
				8'b1001000: c <= 9'b101101;
				8'b111000: c <= 9'b100111110;
				8'b110001: c <= 9'b1101110;
				8'b1010111: c <= 9'b10110011;
				8'b1001110: c <= 9'b110011010;
				8'b1101010: c <= 9'b11;
				8'b1001001: c <= 9'b110011110;
				8'b1100000: c <= 9'b11001011;
				8'b110111: c <= 9'b10111101;
				8'b1011101: c <= 9'b100100101;
				8'b1011011: c <= 9'b1100;
				8'b111001: c <= 9'b10000101;
				8'b1001010: c <= 9'b100101000;
				8'b110011: c <= 9'b100010101;
				8'b1101100: c <= 9'b111110110;
				8'b1110111: c <= 9'b10111111;
				8'b101011: c <= 9'b10101000;
				8'b1101011: c <= 9'b101000110;
				8'b111100: c <= 9'b11000000;
				8'b1000111: c <= 9'b1101000;
				8'b1011111: c <= 9'b11011010;
				8'b1110100: c <= 9'b1111011;
				8'b101101: c <= 9'b100011100;
				8'b1010011: c <= 9'b100100011;
				8'b1100001: c <= 9'b10000000;
				8'b110101: c <= 9'b100101110;
				8'b1000100: c <= 9'b100101001;
				8'b1010001: c <= 9'b10100101;
				8'b1010100: c <= 9'b100000110;
				8'b1100110: c <= 9'b11101101;
				8'b101010: c <= 9'b10001110;
				8'b1011110: c <= 9'b101010100;
				8'b1100111: c <= 9'b11001111;
				8'b1011010: c <= 9'b11000100;
				8'b1000010: c <= 9'b10011101;
				8'b111101: c <= 9'b11010011;
				8'b110000: c <= 9'b100011001;
				8'b111110: c <= 9'b10111011;
				8'b1100010: c <= 9'b10111101;
				8'b1110000: c <= 9'b101111001;
				8'b1101001: c <= 9'b10101;
				8'b1110011: c <= 9'b10111000;
				8'b1001100: c <= 9'b11101;
				8'b100001: c <= 9'b1110010;
				8'b1000110: c <= 9'b11010001;
				8'b1110010: c <= 9'b1000011;
				8'b1010000: c <= 9'b101100100;
				8'b1111010: c <= 9'b100011101;
				8'b1010101: c <= 9'b111100100;
				8'b111011: c <= 9'b101001001;
				8'b1001101: c <= 9'b110111111;
				8'b111111: c <= 9'b110000101;
				8'b1101110: c <= 9'b11101111;
				8'b1111011: c <= 9'b11011011;
				8'b1001011: c <= 9'b100101101;
				8'b1101111: c <= 9'b101000110;
				8'b1101000: c <= 9'b110000110;
				8'b101100: c <= 9'b100001100;
				8'b100100: c <= 9'b100000000;
				8'b1111000: c <= 9'b110100000;
				8'b1000101: c <= 9'b1111100;
				8'b1011001: c <= 9'b100110000;
				8'b110100: c <= 9'b11011000;
				8'b1111001: c <= 9'b111101101;
				8'b1110001: c <= 9'b110100000;
				8'b1001111: c <= 9'b100000011;
				8'b1100101: c <= 9'b10101101;
				8'b1111110: c <= 9'b110001011;
				8'b1111100: c <= 9'b110110011;
				8'b1010110: c <= 9'b101110001;
				8'b110010: c <= 9'b1110010;
				8'b1101101: c <= 9'b111000101;
				8'b100011: c <= 9'b101001111;
				8'b1110101: c <= 9'b110100110;
				8'b1111101: c <= 9'b100010000;
				8'b101001: c <= 9'b10101001;
				8'b1010010: c <= 9'b10001000;
				8'b1011000: c <= 9'b1000001;
				8'b101110: c <= 9'b11110100;
				8'b1000001: c <= 9'b10110110;
				default: c <= 9'b0;
			endcase
			9'b100101010 : case(di)
				8'b1000011: c <= 9'b101101101;
				8'b101000: c <= 9'b11100010;
				8'b111010: c <= 9'b10001011;
				8'b110110: c <= 9'b111011111;
				8'b1100100: c <= 9'b1100;
				8'b1000000: c <= 9'b1011111;
				8'b1110110: c <= 9'b101011000;
				8'b100101: c <= 9'b110011;
				8'b101111: c <= 9'b1001010;
				8'b100110: c <= 9'b100000101;
				8'b1100011: c <= 9'b111110001;
				8'b1001000: c <= 9'b110110011;
				8'b111000: c <= 9'b1101010;
				8'b110001: c <= 9'b100010110;
				8'b1010111: c <= 9'b100010101;
				8'b1001110: c <= 9'b101001011;
				8'b1101010: c <= 9'b10101011;
				8'b1001001: c <= 9'b111100001;
				8'b1100000: c <= 9'b110000111;
				8'b110111: c <= 9'b101110111;
				8'b1011101: c <= 9'b10111001;
				8'b1011011: c <= 9'b11010101;
				8'b111001: c <= 9'b10101;
				8'b1001010: c <= 9'b100001111;
				8'b110011: c <= 9'b111000110;
				8'b1101100: c <= 9'b111100;
				8'b1110111: c <= 9'b11001100;
				8'b101011: c <= 9'b101100110;
				8'b1101011: c <= 9'b111101010;
				8'b111100: c <= 9'b11000011;
				8'b1000111: c <= 9'b110010;
				8'b1011111: c <= 9'b1100110;
				8'b1110100: c <= 9'b101000101;
				8'b101101: c <= 9'b1011;
				8'b1010011: c <= 9'b1000010;
				8'b1100001: c <= 9'b101001111;
				8'b110101: c <= 9'b11110011;
				8'b1000100: c <= 9'b111111111;
				8'b1010001: c <= 9'b11010100;
				8'b1010100: c <= 9'b111100011;
				8'b1100110: c <= 9'b1011110;
				8'b101010: c <= 9'b10000101;
				8'b1011110: c <= 9'b111100101;
				8'b1100111: c <= 9'b10010101;
				8'b1011010: c <= 9'b1010111;
				8'b1000010: c <= 9'b1001011;
				8'b111101: c <= 9'b110011011;
				8'b110000: c <= 9'b1000110;
				8'b111110: c <= 9'b1101100;
				8'b1100010: c <= 9'b111101101;
				8'b1110000: c <= 9'b101001001;
				8'b1101001: c <= 9'b101010010;
				8'b1110011: c <= 9'b101101010;
				8'b1001100: c <= 9'b101001001;
				8'b100001: c <= 9'b1000001;
				8'b1000110: c <= 9'b110011000;
				8'b1110010: c <= 9'b110000111;
				8'b1010000: c <= 9'b110001000;
				8'b1111010: c <= 9'b101001110;
				8'b1010101: c <= 9'b1110000;
				8'b111011: c <= 9'b11100001;
				8'b1001101: c <= 9'b111111000;
				8'b111111: c <= 9'b10000101;
				8'b1101110: c <= 9'b111000100;
				8'b1111011: c <= 9'b11010000;
				8'b1001011: c <= 9'b11011;
				8'b1101111: c <= 9'b10110110;
				8'b1101000: c <= 9'b11001101;
				8'b101100: c <= 9'b100101111;
				8'b100100: c <= 9'b1011111;
				8'b1111000: c <= 9'b100110100;
				8'b1000101: c <= 9'b1011;
				8'b1011001: c <= 9'b1100010;
				8'b110100: c <= 9'b110111111;
				8'b1111001: c <= 9'b101011000;
				8'b1110001: c <= 9'b100110101;
				8'b1001111: c <= 9'b110101111;
				8'b1100101: c <= 9'b11;
				8'b1111110: c <= 9'b1100101;
				8'b1111100: c <= 9'b101010010;
				8'b1010110: c <= 9'b110111001;
				8'b110010: c <= 9'b111011101;
				8'b1101101: c <= 9'b10110001;
				8'b100011: c <= 9'b10010100;
				8'b1110101: c <= 9'b110001110;
				8'b1111101: c <= 9'b111111111;
				8'b101001: c <= 9'b10010111;
				8'b1010010: c <= 9'b100001;
				8'b1011000: c <= 9'b101001000;
				8'b101110: c <= 9'b110010011;
				8'b1000001: c <= 9'b101110;
				default: c <= 9'b0;
			endcase
			9'b11010101 : case(di)
				8'b1000011: c <= 9'b101010110;
				8'b101000: c <= 9'b100111000;
				8'b111010: c <= 9'b1110111;
				8'b110110: c <= 9'b1111111;
				8'b1100100: c <= 9'b101110111;
				8'b1000000: c <= 9'b101011110;
				8'b1110110: c <= 9'b11001000;
				8'b100101: c <= 9'b10001010;
				8'b101111: c <= 9'b110011011;
				8'b100110: c <= 9'b101110111;
				8'b1100011: c <= 9'b111010110;
				8'b1001000: c <= 9'b110111001;
				8'b111000: c <= 9'b1111100;
				8'b110001: c <= 9'b101010000;
				8'b1010111: c <= 9'b10101001;
				8'b1001110: c <= 9'b110011100;
				8'b1101010: c <= 9'b11111110;
				8'b1001001: c <= 9'b11101000;
				8'b1100000: c <= 9'b111110110;
				8'b110111: c <= 9'b10101000;
				8'b1011101: c <= 9'b1101000;
				8'b1011011: c <= 9'b110110110;
				8'b111001: c <= 9'b10001001;
				8'b1001010: c <= 9'b110011010;
				8'b110011: c <= 9'b101000111;
				8'b1101100: c <= 9'b100000001;
				8'b1110111: c <= 9'b101001;
				8'b101011: c <= 9'b11101001;
				8'b1101011: c <= 9'b1110000;
				8'b111100: c <= 9'b110011;
				8'b1000111: c <= 9'b11010001;
				8'b1011111: c <= 9'b100010101;
				8'b1110100: c <= 9'b10000110;
				8'b101101: c <= 9'b100010101;
				8'b1010011: c <= 9'b10000;
				8'b1100001: c <= 9'b101000101;
				8'b110101: c <= 9'b101100110;
				8'b1000100: c <= 9'b1001000;
				8'b1010001: c <= 9'b101001010;
				8'b1010100: c <= 9'b10011111;
				8'b1100110: c <= 9'b11010101;
				8'b101010: c <= 9'b1111111;
				8'b1011110: c <= 9'b101111000;
				8'b1100111: c <= 9'b1010101;
				8'b1011010: c <= 9'b10111000;
				8'b1000010: c <= 9'b110101110;
				8'b111101: c <= 9'b111111011;
				8'b110000: c <= 9'b100101101;
				8'b111110: c <= 9'b11110110;
				8'b1100010: c <= 9'b11100001;
				8'b1110000: c <= 9'b111100111;
				8'b1101001: c <= 9'b10000110;
				8'b1110011: c <= 9'b1011011;
				8'b1001100: c <= 9'b111000110;
				8'b100001: c <= 9'b1100101;
				8'b1000110: c <= 9'b111111;
				8'b1110010: c <= 9'b101101110;
				8'b1010000: c <= 9'b111000100;
				8'b1111010: c <= 9'b100101001;
				8'b1010101: c <= 9'b100111001;
				8'b111011: c <= 9'b100010111;
				8'b1001101: c <= 9'b111011010;
				8'b111111: c <= 9'b110100010;
				8'b1101110: c <= 9'b110100001;
				8'b1111011: c <= 9'b10101100;
				8'b1001011: c <= 9'b101001001;
				8'b1101111: c <= 9'b111100001;
				8'b1101000: c <= 9'b111000111;
				8'b101100: c <= 9'b111101111;
				8'b100100: c <= 9'b100001110;
				8'b1111000: c <= 9'b1001111;
				8'b1000101: c <= 9'b101010011;
				8'b1011001: c <= 9'b110101111;
				8'b110100: c <= 9'b111100101;
				8'b1111001: c <= 9'b10110011;
				8'b1110001: c <= 9'b111000100;
				8'b1001111: c <= 9'b11010010;
				8'b1100101: c <= 9'b10001000;
				8'b1111110: c <= 9'b1010011;
				8'b1111100: c <= 9'b10010;
				8'b1010110: c <= 9'b101000110;
				8'b110010: c <= 9'b10010110;
				8'b1101101: c <= 9'b111101101;
				8'b100011: c <= 9'b101001111;
				8'b1110101: c <= 9'b101101100;
				8'b1111101: c <= 9'b101100011;
				8'b101001: c <= 9'b100100101;
				8'b1010010: c <= 9'b110110110;
				8'b1011000: c <= 9'b11010011;
				8'b101110: c <= 9'b10101010;
				8'b1000001: c <= 9'b101001011;
				default: c <= 9'b0;
			endcase
			9'b111100111 : case(di)
				8'b1000011: c <= 9'b101101110;
				8'b101000: c <= 9'b1111000;
				8'b111010: c <= 9'b111101000;
				8'b110110: c <= 9'b110111111;
				8'b1100100: c <= 9'b10011011;
				8'b1000000: c <= 9'b100111011;
				8'b1110110: c <= 9'b110000011;
				8'b100101: c <= 9'b11111011;
				8'b101111: c <= 9'b111100011;
				8'b100110: c <= 9'b111101;
				8'b1100011: c <= 9'b10110101;
				8'b1001000: c <= 9'b101110000;
				8'b111000: c <= 9'b1010101;
				8'b110001: c <= 9'b111010100;
				8'b1010111: c <= 9'b11111011;
				8'b1001110: c <= 9'b100100111;
				8'b1101010: c <= 9'b101011;
				8'b1001001: c <= 9'b100110011;
				8'b1100000: c <= 9'b101110001;
				8'b110111: c <= 9'b101001001;
				8'b1011101: c <= 9'b10011111;
				8'b1011011: c <= 9'b101101010;
				8'b111001: c <= 9'b111110000;
				8'b1001010: c <= 9'b101000001;
				8'b110011: c <= 9'b10001010;
				8'b1101100: c <= 9'b101101111;
				8'b1110111: c <= 9'b10000001;
				8'b101011: c <= 9'b10011111;
				8'b1101011: c <= 9'b110001001;
				8'b111100: c <= 9'b100001;
				8'b1000111: c <= 9'b1101100;
				8'b1011111: c <= 9'b111100011;
				8'b1110100: c <= 9'b100010110;
				8'b101101: c <= 9'b11000111;
				8'b1010011: c <= 9'b11010111;
				8'b1100001: c <= 9'b10111100;
				8'b110101: c <= 9'b11001100;
				8'b1000100: c <= 9'b100100;
				8'b1010001: c <= 9'b10110111;
				8'b1010100: c <= 9'b10010011;
				8'b1100110: c <= 9'b11001011;
				8'b101010: c <= 9'b11100111;
				8'b1011110: c <= 9'b1001;
				8'b1100111: c <= 9'b101101100;
				8'b1011010: c <= 9'b11110010;
				8'b1000010: c <= 9'b11101100;
				8'b111101: c <= 9'b1111001;
				8'b110000: c <= 9'b10110010;
				8'b111110: c <= 9'b110111111;
				8'b1100010: c <= 9'b1011110;
				8'b1110000: c <= 9'b1000000;
				8'b1101001: c <= 9'b110110;
				8'b1110011: c <= 9'b11111;
				8'b1001100: c <= 9'b111000101;
				8'b100001: c <= 9'b1000011;
				8'b1000110: c <= 9'b10010001;
				8'b1110010: c <= 9'b11011;
				8'b1010000: c <= 9'b10001001;
				8'b1111010: c <= 9'b111110101;
				8'b1010101: c <= 9'b100111101;
				8'b111011: c <= 9'b101111000;
				8'b1001101: c <= 9'b101;
				8'b111111: c <= 9'b10001110;
				8'b1101110: c <= 9'b1011100;
				8'b1111011: c <= 9'b111011101;
				8'b1001011: c <= 9'b110110010;
				8'b1101111: c <= 9'b111101010;
				8'b1101000: c <= 9'b10011111;
				8'b101100: c <= 9'b101101000;
				8'b100100: c <= 9'b101101101;
				8'b1111000: c <= 9'b1010110;
				8'b1000101: c <= 9'b1100111;
				8'b1011001: c <= 9'b100110;
				8'b110100: c <= 9'b111100000;
				8'b1111001: c <= 9'b110110111;
				8'b1110001: c <= 9'b101110110;
				8'b1001111: c <= 9'b11110110;
				8'b1100101: c <= 9'b100;
				8'b1111110: c <= 9'b101000111;
				8'b1111100: c <= 9'b110001110;
				8'b1010110: c <= 9'b10110010;
				8'b110010: c <= 9'b10011111;
				8'b1101101: c <= 9'b101000010;
				8'b100011: c <= 9'b101100100;
				8'b1110101: c <= 9'b110011100;
				8'b1111101: c <= 9'b100100000;
				8'b101001: c <= 9'b101000110;
				8'b1010010: c <= 9'b10110100;
				8'b1011000: c <= 9'b110111000;
				8'b101110: c <= 9'b111010001;
				8'b1000001: c <= 9'b111010100;
				default: c <= 9'b0;
			endcase
			9'b100110011 : case(di)
				8'b1000011: c <= 9'b10100;
				8'b101000: c <= 9'b1110011;
				8'b111010: c <= 9'b1110111;
				8'b110110: c <= 9'b10010100;
				8'b1100100: c <= 9'b10011001;
				8'b1000000: c <= 9'b10101010;
				8'b1110110: c <= 9'b1101100;
				8'b100101: c <= 9'b10110010;
				8'b101111: c <= 9'b10101011;
				8'b100110: c <= 9'b10000110;
				8'b1100011: c <= 9'b1110011;
				8'b1001000: c <= 9'b10010111;
				8'b111000: c <= 9'b11001010;
				8'b110001: c <= 9'b10011111;
				8'b1010111: c <= 9'b100011100;
				8'b1001110: c <= 9'b101110000;
				8'b1101010: c <= 9'b10011001;
				8'b1001001: c <= 9'b111100110;
				8'b1100000: c <= 9'b100111110;
				8'b110111: c <= 9'b11110111;
				8'b1011101: c <= 9'b1010011;
				8'b1011011: c <= 9'b110110010;
				8'b111001: c <= 9'b11011101;
				8'b1001010: c <= 9'b1100100;
				8'b110011: c <= 9'b1111000;
				8'b1101100: c <= 9'b10100010;
				8'b1110111: c <= 9'b10100000;
				8'b101011: c <= 9'b110100001;
				8'b1101011: c <= 9'b100001110;
				8'b111100: c <= 9'b11010001;
				8'b1000111: c <= 9'b101011000;
				8'b1011111: c <= 9'b10010000;
				8'b1110100: c <= 9'b100101000;
				8'b101101: c <= 9'b10001011;
				8'b1010011: c <= 9'b110101001;
				8'b1100001: c <= 9'b1001011;
				8'b110101: c <= 9'b101110110;
				8'b1000100: c <= 9'b111010100;
				8'b1010001: c <= 9'b11110001;
				8'b1010100: c <= 9'b11110010;
				8'b1100110: c <= 9'b100011000;
				8'b101010: c <= 9'b10111101;
				8'b1011110: c <= 9'b10111011;
				8'b1100111: c <= 9'b1100110;
				8'b1011010: c <= 9'b111101111;
				8'b1000010: c <= 9'b101100011;
				8'b111101: c <= 9'b101001111;
				8'b110000: c <= 9'b110100010;
				8'b111110: c <= 9'b101001010;
				8'b1100010: c <= 9'b1110001;
				8'b1110000: c <= 9'b10001100;
				8'b1101001: c <= 9'b101000110;
				8'b1110011: c <= 9'b100000010;
				8'b1001100: c <= 9'b110001111;
				8'b100001: c <= 9'b1101101;
				8'b1000110: c <= 9'b110111100;
				8'b1110010: c <= 9'b10001011;
				8'b1010000: c <= 9'b11111000;
				8'b1111010: c <= 9'b101010110;
				8'b1010101: c <= 9'b11001001;
				8'b111011: c <= 9'b100000110;
				8'b1001101: c <= 9'b100101;
				8'b111111: c <= 9'b101101010;
				8'b1101110: c <= 9'b100011101;
				8'b1111011: c <= 9'b100011111;
				8'b1001011: c <= 9'b101110111;
				8'b1101111: c <= 9'b1;
				8'b1101000: c <= 9'b1011111;
				8'b101100: c <= 9'b11011000;
				8'b100100: c <= 9'b101100111;
				8'b1111000: c <= 9'b1101100;
				8'b1000101: c <= 9'b110011111;
				8'b1011001: c <= 9'b11100011;
				8'b110100: c <= 9'b100001100;
				8'b1111001: c <= 9'b110011000;
				8'b1110001: c <= 9'b101110000;
				8'b1001111: c <= 9'b111011101;
				8'b1100101: c <= 9'b110101001;
				8'b1111110: c <= 9'b111111000;
				8'b1111100: c <= 9'b110001011;
				8'b1010110: c <= 9'b10100101;
				8'b110010: c <= 9'b101100010;
				8'b1101101: c <= 9'b101101001;
				8'b100011: c <= 9'b100000100;
				8'b1110101: c <= 9'b101100001;
				8'b1111101: c <= 9'b11100000;
				8'b101001: c <= 9'b10;
				8'b1010010: c <= 9'b10001011;
				8'b1011000: c <= 9'b100011000;
				8'b101110: c <= 9'b111001;
				8'b1000001: c <= 9'b100001111;
				default: c <= 9'b0;
			endcase
			9'b11001001 : case(di)
				8'b1000011: c <= 9'b100010011;
				8'b101000: c <= 9'b111010000;
				8'b111010: c <= 9'b110000001;
				8'b110110: c <= 9'b100111111;
				8'b1100100: c <= 9'b1000011;
				8'b1000000: c <= 9'b10001010;
				8'b1110110: c <= 9'b1011010;
				8'b100101: c <= 9'b110101010;
				8'b101111: c <= 9'b110110110;
				8'b100110: c <= 9'b1100111;
				8'b1100011: c <= 9'b110111001;
				8'b1001000: c <= 9'b100100111;
				8'b111000: c <= 9'b100010101;
				8'b110001: c <= 9'b100111001;
				8'b1010111: c <= 9'b1100001;
				8'b1001110: c <= 9'b101100100;
				8'b1101010: c <= 9'b100;
				8'b1001001: c <= 9'b11011100;
				8'b1100000: c <= 9'b10100011;
				8'b110111: c <= 9'b1100100;
				8'b1011101: c <= 9'b11010;
				8'b1011011: c <= 9'b101010;
				8'b111001: c <= 9'b1101110;
				8'b1001010: c <= 9'b11101000;
				8'b110011: c <= 9'b11011101;
				8'b1101100: c <= 9'b10100011;
				8'b1110111: c <= 9'b1100010;
				8'b101011: c <= 9'b11000111;
				8'b1101011: c <= 9'b11010011;
				8'b111100: c <= 9'b1001101;
				8'b1000111: c <= 9'b11111101;
				8'b1011111: c <= 9'b11010001;
				8'b1110100: c <= 9'b11001010;
				8'b101101: c <= 9'b1111001;
				8'b1010011: c <= 9'b10110110;
				8'b1100001: c <= 9'b101011001;
				8'b110101: c <= 9'b111111010;
				8'b1000100: c <= 9'b1001010;
				8'b1010001: c <= 9'b100101000;
				8'b1010100: c <= 9'b111110110;
				8'b1100110: c <= 9'b100010010;
				8'b101010: c <= 9'b11000010;
				8'b1011110: c <= 9'b101111001;
				8'b1100111: c <= 9'b10010001;
				8'b1011010: c <= 9'b1010110;
				8'b1000010: c <= 9'b101000111;
				8'b111101: c <= 9'b110;
				8'b110000: c <= 9'b1100101;
				8'b111110: c <= 9'b10110111;
				8'b1100010: c <= 9'b11100111;
				8'b1110000: c <= 9'b11001101;
				8'b1101001: c <= 9'b11100011;
				8'b1110011: c <= 9'b110101;
				8'b1001100: c <= 9'b100100101;
				8'b100001: c <= 9'b100001110;
				8'b1000110: c <= 9'b100101011;
				8'b1110010: c <= 9'b110101;
				8'b1010000: c <= 9'b110010010;
				8'b1111010: c <= 9'b10110011;
				8'b1010101: c <= 9'b11101100;
				8'b111011: c <= 9'b110010101;
				8'b1001101: c <= 9'b100001100;
				8'b111111: c <= 9'b100000011;
				8'b1101110: c <= 9'b110000010;
				8'b1111011: c <= 9'b101111001;
				8'b1001011: c <= 9'b101101010;
				8'b1101111: c <= 9'b100001011;
				8'b1101000: c <= 9'b1001101;
				8'b101100: c <= 9'b110100110;
				8'b100100: c <= 9'b11111110;
				8'b1111000: c <= 9'b100010010;
				8'b1000101: c <= 9'b11001011;
				8'b1011001: c <= 9'b111000011;
				8'b110100: c <= 9'b101001010;
				8'b1111001: c <= 9'b100110110;
				8'b1110001: c <= 9'b101101000;
				8'b1001111: c <= 9'b1;
				8'b1100101: c <= 9'b1111101;
				8'b1111110: c <= 9'b111100011;
				8'b1111100: c <= 9'b110101001;
				8'b1010110: c <= 9'b10101100;
				8'b110010: c <= 9'b111001110;
				8'b1101101: c <= 9'b101011000;
				8'b100011: c <= 9'b111010110;
				8'b1110101: c <= 9'b101011001;
				8'b1111101: c <= 9'b110100;
				8'b101001: c <= 9'b10110110;
				8'b1010010: c <= 9'b110001011;
				8'b1011000: c <= 9'b10000011;
				8'b101110: c <= 9'b110100111;
				8'b1000001: c <= 9'b10000010;
				default: c <= 9'b0;
			endcase
			9'b101100010 : case(di)
				8'b1000011: c <= 9'b101001100;
				8'b101000: c <= 9'b11000000;
				8'b111010: c <= 9'b100101010;
				8'b110110: c <= 9'b101011001;
				8'b1100100: c <= 9'b10000101;
				8'b1000000: c <= 9'b111000110;
				8'b1110110: c <= 9'b110000001;
				8'b100101: c <= 9'b10101;
				8'b101111: c <= 9'b1110100;
				8'b100110: c <= 9'b100010011;
				8'b1100011: c <= 9'b101000001;
				8'b1001000: c <= 9'b101100000;
				8'b111000: c <= 9'b110011011;
				8'b110001: c <= 9'b100111010;
				8'b1010111: c <= 9'b110100111;
				8'b1001110: c <= 9'b101011000;
				8'b1101010: c <= 9'b101100010;
				8'b1001001: c <= 9'b10110111;
				8'b1100000: c <= 9'b110000101;
				8'b110111: c <= 9'b100010000;
				8'b1011101: c <= 9'b11101001;
				8'b1011011: c <= 9'b10011001;
				8'b111001: c <= 9'b101000101;
				8'b1001010: c <= 9'b1111011;
				8'b110011: c <= 9'b111111111;
				8'b1101100: c <= 9'b1010010;
				8'b1110111: c <= 9'b110111011;
				8'b101011: c <= 9'b1010110;
				8'b1101011: c <= 9'b1110101;
				8'b111100: c <= 9'b110001000;
				8'b1000111: c <= 9'b100001110;
				8'b1011111: c <= 9'b110000110;
				8'b1110100: c <= 9'b1010101;
				8'b101101: c <= 9'b100101001;
				8'b1010011: c <= 9'b100010111;
				8'b1100001: c <= 9'b1;
				8'b110101: c <= 9'b111000111;
				8'b1000100: c <= 9'b111011011;
				8'b1010001: c <= 9'b110111;
				8'b1010100: c <= 9'b110010100;
				8'b1100110: c <= 9'b110001101;
				8'b101010: c <= 9'b110000011;
				8'b1011110: c <= 9'b11100110;
				8'b1100111: c <= 9'b1100111;
				8'b1011010: c <= 9'b1011110;
				8'b1000010: c <= 9'b1101001;
				8'b111101: c <= 9'b110000110;
				8'b110000: c <= 9'b100011100;
				8'b111110: c <= 9'b110011100;
				8'b1100010: c <= 9'b1011011;
				8'b1110000: c <= 9'b110000010;
				8'b1101001: c <= 9'b11011010;
				8'b1110011: c <= 9'b11101;
				8'b1001100: c <= 9'b100101100;
				8'b100001: c <= 9'b111000110;
				8'b1000110: c <= 9'b111101111;
				8'b1110010: c <= 9'b1000;
				8'b1010000: c <= 9'b100010100;
				8'b1111010: c <= 9'b101001110;
				8'b1010101: c <= 9'b110010101;
				8'b111011: c <= 9'b10;
				8'b1001101: c <= 9'b110101010;
				8'b111111: c <= 9'b110100111;
				8'b1101110: c <= 9'b10100011;
				8'b1111011: c <= 9'b110001111;
				8'b1001011: c <= 9'b10101101;
				8'b1101111: c <= 9'b100110110;
				8'b1101000: c <= 9'b1010001;
				8'b101100: c <= 9'b1001;
				8'b100100: c <= 9'b10011100;
				8'b1111000: c <= 9'b111001101;
				8'b1000101: c <= 9'b11000100;
				8'b1011001: c <= 9'b11101;
				8'b110100: c <= 9'b1011110;
				8'b1111001: c <= 9'b11011110;
				8'b1110001: c <= 9'b11000;
				8'b1001111: c <= 9'b1110101;
				8'b1100101: c <= 9'b1111101;
				8'b1111110: c <= 9'b100010;
				8'b1111100: c <= 9'b101110;
				8'b1010110: c <= 9'b10110101;
				8'b110010: c <= 9'b11011100;
				8'b1101101: c <= 9'b11000010;
				8'b100011: c <= 9'b111010000;
				8'b1110101: c <= 9'b10001111;
				8'b1111101: c <= 9'b110011011;
				8'b101001: c <= 9'b101110111;
				8'b1010010: c <= 9'b1011011;
				8'b1011000: c <= 9'b11110;
				8'b101110: c <= 9'b110000101;
				8'b1000001: c <= 9'b110100;
				default: c <= 9'b0;
			endcase
			9'b1001000 : case(di)
				8'b1000011: c <= 9'b1010010;
				8'b101000: c <= 9'b101110001;
				8'b111010: c <= 9'b11100101;
				8'b110110: c <= 9'b110110;
				8'b1100100: c <= 9'b111110000;
				8'b1000000: c <= 9'b110001101;
				8'b1110110: c <= 9'b100101100;
				8'b100101: c <= 9'b100100000;
				8'b101111: c <= 9'b100100000;
				8'b100110: c <= 9'b111001000;
				8'b1100011: c <= 9'b100100011;
				8'b1001000: c <= 9'b101100101;
				8'b111000: c <= 9'b10110010;
				8'b110001: c <= 9'b100111010;
				8'b1010111: c <= 9'b10100111;
				8'b1001110: c <= 9'b100001110;
				8'b1101010: c <= 9'b11110001;
				8'b1001001: c <= 9'b110111100;
				8'b1100000: c <= 9'b1110011;
				8'b110111: c <= 9'b101000;
				8'b1011101: c <= 9'b101101010;
				8'b1011011: c <= 9'b1001000;
				8'b111001: c <= 9'b101000111;
				8'b1001010: c <= 9'b100010101;
				8'b110011: c <= 9'b111011010;
				8'b1101100: c <= 9'b111100111;
				8'b1110111: c <= 9'b100111101;
				8'b101011: c <= 9'b110010011;
				8'b1101011: c <= 9'b101101011;
				8'b111100: c <= 9'b110101101;
				8'b1000111: c <= 9'b10010011;
				8'b1011111: c <= 9'b10100010;
				8'b1110100: c <= 9'b110010011;
				8'b101101: c <= 9'b100101110;
				8'b1010011: c <= 9'b11100110;
				8'b1100001: c <= 9'b11010010;
				8'b110101: c <= 9'b111011010;
				8'b1000100: c <= 9'b101100;
				8'b1010001: c <= 9'b10111011;
				8'b1010100: c <= 9'b10110111;
				8'b1100110: c <= 9'b110100101;
				8'b101010: c <= 9'b10000011;
				8'b1011110: c <= 9'b110011000;
				8'b1100111: c <= 9'b111011111;
				8'b1011010: c <= 9'b10001010;
				8'b1000010: c <= 9'b110001000;
				8'b111101: c <= 9'b100110000;
				8'b110000: c <= 9'b100100111;
				8'b111110: c <= 9'b111101100;
				8'b1100010: c <= 9'b110100;
				8'b1110000: c <= 9'b110100001;
				8'b1101001: c <= 9'b1111011;
				8'b1110011: c <= 9'b110100011;
				8'b1001100: c <= 9'b101000100;
				8'b100001: c <= 9'b10111010;
				8'b1000110: c <= 9'b10011101;
				8'b1110010: c <= 9'b101011110;
				8'b1010000: c <= 9'b101100101;
				8'b1111010: c <= 9'b101010001;
				8'b1010101: c <= 9'b100000111;
				8'b111011: c <= 9'b110000011;
				8'b1001101: c <= 9'b101001110;
				8'b111111: c <= 9'b111001101;
				8'b1101110: c <= 9'b101110111;
				8'b1111011: c <= 9'b10100;
				8'b1001011: c <= 9'b11110011;
				8'b1101111: c <= 9'b10100000;
				8'b1101000: c <= 9'b110011100;
				8'b101100: c <= 9'b101101001;
				8'b100100: c <= 9'b11111110;
				8'b1111000: c <= 9'b111110110;
				8'b1000101: c <= 9'b100001001;
				8'b1011001: c <= 9'b11000;
				8'b110100: c <= 9'b11101011;
				8'b1111001: c <= 9'b101110011;
				8'b1110001: c <= 9'b10001111;
				8'b1001111: c <= 9'b110110100;
				8'b1100101: c <= 9'b101010;
				8'b1111110: c <= 9'b111010100;
				8'b1111100: c <= 9'b10101011;
				8'b1010110: c <= 9'b1011010;
				8'b110010: c <= 9'b10110011;
				8'b1101101: c <= 9'b1010110;
				8'b100011: c <= 9'b110110100;
				8'b1110101: c <= 9'b101110001;
				8'b1111101: c <= 9'b1000001;
				8'b101001: c <= 9'b11010101;
				8'b1010010: c <= 9'b101101111;
				8'b1011000: c <= 9'b110100110;
				8'b101110: c <= 9'b100001110;
				8'b1000001: c <= 9'b10001000;
				default: c <= 9'b0;
			endcase
			9'b111010010 : case(di)
				8'b1000011: c <= 9'b100110;
				8'b101000: c <= 9'b100000011;
				8'b111010: c <= 9'b110101110;
				8'b110110: c <= 9'b1101110;
				8'b1100100: c <= 9'b11111011;
				8'b1000000: c <= 9'b10101110;
				8'b1110110: c <= 9'b111101100;
				8'b100101: c <= 9'b11111100;
				8'b101111: c <= 9'b11011010;
				8'b100110: c <= 9'b101101000;
				8'b1100011: c <= 9'b100011011;
				8'b1001000: c <= 9'b10101101;
				8'b111000: c <= 9'b11110;
				8'b110001: c <= 9'b110101001;
				8'b1010111: c <= 9'b100101100;
				8'b1001110: c <= 9'b10011010;
				8'b1101010: c <= 9'b1001011;
				8'b1001001: c <= 9'b10110001;
				8'b1100000: c <= 9'b10011011;
				8'b110111: c <= 9'b101011010;
				8'b1011101: c <= 9'b111100100;
				8'b1011011: c <= 9'b10110101;
				8'b111001: c <= 9'b111001010;
				8'b1001010: c <= 9'b100100110;
				8'b110011: c <= 9'b110111110;
				8'b1101100: c <= 9'b10101111;
				8'b1110111: c <= 9'b100101010;
				8'b101011: c <= 9'b1111010;
				8'b1101011: c <= 9'b10011;
				8'b111100: c <= 9'b10100;
				8'b1000111: c <= 9'b100100110;
				8'b1011111: c <= 9'b100000111;
				8'b1110100: c <= 9'b11100011;
				8'b101101: c <= 9'b10101000;
				8'b1010011: c <= 9'b100011001;
				8'b1100001: c <= 9'b10000000;
				8'b110101: c <= 9'b101001110;
				8'b1000100: c <= 9'b101011110;
				8'b1010001: c <= 9'b11101001;
				8'b1010100: c <= 9'b1101001;
				8'b1100110: c <= 9'b110110000;
				8'b101010: c <= 9'b11100011;
				8'b1011110: c <= 9'b110000001;
				8'b1100111: c <= 9'b11100010;
				8'b1011010: c <= 9'b111011;
				8'b1000010: c <= 9'b111101001;
				8'b111101: c <= 9'b110010;
				8'b110000: c <= 9'b110101100;
				8'b111110: c <= 9'b11100;
				8'b1100010: c <= 9'b1011011;
				8'b1110000: c <= 9'b11001;
				8'b1101001: c <= 9'b110010;
				8'b1110011: c <= 9'b100011001;
				8'b1001100: c <= 9'b100010101;
				8'b100001: c <= 9'b1100100;
				8'b1000110: c <= 9'b10101111;
				8'b1110010: c <= 9'b10001011;
				8'b1010000: c <= 9'b100111110;
				8'b1111010: c <= 9'b10100000;
				8'b1010101: c <= 9'b100111001;
				8'b111011: c <= 9'b100110011;
				8'b1001101: c <= 9'b101011011;
				8'b111111: c <= 9'b10000101;
				8'b1101110: c <= 9'b100000100;
				8'b1111011: c <= 9'b100110110;
				8'b1001011: c <= 9'b100010111;
				8'b1101111: c <= 9'b100101100;
				8'b1101000: c <= 9'b10111000;
				8'b101100: c <= 9'b111000110;
				8'b100100: c <= 9'b11001001;
				8'b1111000: c <= 9'b1110100;
				8'b1000101: c <= 9'b100011000;
				8'b1011001: c <= 9'b1110001;
				8'b110100: c <= 9'b110100010;
				8'b1111001: c <= 9'b111001;
				8'b1110001: c <= 9'b110000101;
				8'b1001111: c <= 9'b100000011;
				8'b1100101: c <= 9'b111011111;
				8'b1111110: c <= 9'b10100000;
				8'b1111100: c <= 9'b10001101;
				8'b1010110: c <= 9'b111101111;
				8'b110010: c <= 9'b110000010;
				8'b1101101: c <= 9'b100011111;
				8'b100011: c <= 9'b101000;
				8'b1110101: c <= 9'b1100000;
				8'b1111101: c <= 9'b10110;
				8'b101001: c <= 9'b101110001;
				8'b1010010: c <= 9'b111011100;
				8'b1011000: c <= 9'b10110111;
				8'b101110: c <= 9'b110110111;
				8'b1000001: c <= 9'b110110;
				default: c <= 9'b0;
			endcase
			9'b111001000 : case(di)
				8'b1000011: c <= 9'b101;
				8'b101000: c <= 9'b100010010;
				8'b111010: c <= 9'b101000111;
				8'b110110: c <= 9'b1100;
				8'b1100100: c <= 9'b100110000;
				8'b1000000: c <= 9'b11101000;
				8'b1110110: c <= 9'b110101100;
				8'b100101: c <= 9'b1011001;
				8'b101111: c <= 9'b111001101;
				8'b100110: c <= 9'b100101101;
				8'b1100011: c <= 9'b110000110;
				8'b1001000: c <= 9'b11110101;
				8'b111000: c <= 9'b11001101;
				8'b110001: c <= 9'b101011010;
				8'b1010111: c <= 9'b111011010;
				8'b1001110: c <= 9'b100101010;
				8'b1101010: c <= 9'b1101001;
				8'b1001001: c <= 9'b10101;
				8'b1100000: c <= 9'b100100101;
				8'b110111: c <= 9'b10101100;
				8'b1011101: c <= 9'b11011001;
				8'b1011011: c <= 9'b111000111;
				8'b111001: c <= 9'b110111110;
				8'b1001010: c <= 9'b11010;
				8'b110011: c <= 9'b1100;
				8'b1101100: c <= 9'b10011000;
				8'b1110111: c <= 9'b1010010;
				8'b101011: c <= 9'b101000110;
				8'b1101011: c <= 9'b10100011;
				8'b111100: c <= 9'b11111;
				8'b1000111: c <= 9'b111111110;
				8'b1011111: c <= 9'b101000100;
				8'b1110100: c <= 9'b1010110;
				8'b101101: c <= 9'b11011011;
				8'b1010011: c <= 9'b111010100;
				8'b1100001: c <= 9'b1100111;
				8'b110101: c <= 9'b101000;
				8'b1000100: c <= 9'b110011100;
				8'b1010001: c <= 9'b101111110;
				8'b1010100: c <= 9'b10100100;
				8'b1100110: c <= 9'b1001110;
				8'b101010: c <= 9'b11110;
				8'b1011110: c <= 9'b111011111;
				8'b1100111: c <= 9'b1011100;
				8'b1011010: c <= 9'b1110101;
				8'b1000010: c <= 9'b101010001;
				8'b111101: c <= 9'b10110;
				8'b110000: c <= 9'b1000111;
				8'b111110: c <= 9'b111010;
				8'b1100010: c <= 9'b110001;
				8'b1110000: c <= 9'b110110110;
				8'b1101001: c <= 9'b110010101;
				8'b1110011: c <= 9'b101011;
				8'b1001100: c <= 9'b10110011;
				8'b100001: c <= 9'b11101111;
				8'b1000110: c <= 9'b110001111;
				8'b1110010: c <= 9'b100011111;
				8'b1010000: c <= 9'b10100000;
				8'b1111010: c <= 9'b1110011;
				8'b1010101: c <= 9'b111011011;
				8'b111011: c <= 9'b10111101;
				8'b1001101: c <= 9'b111000111;
				8'b111111: c <= 9'b111101001;
				8'b1101110: c <= 9'b100100010;
				8'b1111011: c <= 9'b10101110;
				8'b1001011: c <= 9'b10111010;
				8'b1101111: c <= 9'b101001011;
				8'b1101000: c <= 9'b11110;
				8'b101100: c <= 9'b111111001;
				8'b100100: c <= 9'b111001111;
				8'b1111000: c <= 9'b111010;
				8'b1000101: c <= 9'b10000;
				8'b1011001: c <= 9'b1001110;
				8'b110100: c <= 9'b101011;
				8'b1111001: c <= 9'b110101010;
				8'b1110001: c <= 9'b100110100;
				8'b1001111: c <= 9'b10011101;
				8'b1100101: c <= 9'b111011111;
				8'b1111110: c <= 9'b100110010;
				8'b1111100: c <= 9'b110011110;
				8'b1010110: c <= 9'b1000001;
				8'b110010: c <= 9'b11110100;
				8'b1101101: c <= 9'b111111;
				8'b100011: c <= 9'b101001111;
				8'b1110101: c <= 9'b100100001;
				8'b1111101: c <= 9'b100100000;
				8'b101001: c <= 9'b111101;
				8'b1010010: c <= 9'b110001101;
				8'b1011000: c <= 9'b101010101;
				8'b101110: c <= 9'b101111110;
				8'b1000001: c <= 9'b10001111;
				default: c <= 9'b0;
			endcase
			9'b10011111 : case(di)
				8'b1000011: c <= 9'b111110011;
				8'b101000: c <= 9'b1101;
				8'b111010: c <= 9'b111001100;
				8'b110110: c <= 9'b1101111;
				8'b1100100: c <= 9'b111000;
				8'b1000000: c <= 9'b10111010;
				8'b1110110: c <= 9'b1011001;
				8'b100101: c <= 9'b111110001;
				8'b101111: c <= 9'b111110000;
				8'b100110: c <= 9'b111001001;
				8'b1100011: c <= 9'b111000010;
				8'b1001000: c <= 9'b101101;
				8'b111000: c <= 9'b101101011;
				8'b110001: c <= 9'b111010010;
				8'b1010111: c <= 9'b100101000;
				8'b1001110: c <= 9'b11001010;
				8'b1101010: c <= 9'b10010000;
				8'b1001001: c <= 9'b11000001;
				8'b1100000: c <= 9'b1100100;
				8'b110111: c <= 9'b110100010;
				8'b1011101: c <= 9'b111101010;
				8'b1011011: c <= 9'b10101100;
				8'b111001: c <= 9'b110010110;
				8'b1001010: c <= 9'b11001100;
				8'b110011: c <= 9'b100100010;
				8'b1101100: c <= 9'b110011110;
				8'b1110111: c <= 9'b111010111;
				8'b101011: c <= 9'b110110101;
				8'b1101011: c <= 9'b1111110;
				8'b111100: c <= 9'b110011110;
				8'b1000111: c <= 9'b1100000;
				8'b1011111: c <= 9'b111110101;
				8'b1110100: c <= 9'b11110111;
				8'b101101: c <= 9'b1010101;
				8'b1010011: c <= 9'b10111;
				8'b1100001: c <= 9'b111001010;
				8'b110101: c <= 9'b11100001;
				8'b1000100: c <= 9'b100010101;
				8'b1010001: c <= 9'b110011011;
				8'b1010100: c <= 9'b1111100;
				8'b1100110: c <= 9'b11101111;
				8'b101010: c <= 9'b100010011;
				8'b1011110: c <= 9'b11110100;
				8'b1100111: c <= 9'b10110011;
				8'b1011010: c <= 9'b110111100;
				8'b1000010: c <= 9'b1000010;
				8'b111101: c <= 9'b10111111;
				8'b110000: c <= 9'b10001111;
				8'b111110: c <= 9'b11001101;
				8'b1100010: c <= 9'b100;
				8'b1110000: c <= 9'b11001001;
				8'b1101001: c <= 9'b100100010;
				8'b1110011: c <= 9'b11000100;
				8'b1001100: c <= 9'b1101010;
				8'b100001: c <= 9'b111010001;
				8'b1000110: c <= 9'b11101000;
				8'b1110010: c <= 9'b101001111;
				8'b1010000: c <= 9'b10110001;
				8'b1111010: c <= 9'b111101000;
				8'b1010101: c <= 9'b1000100;
				8'b111011: c <= 9'b100010001;
				8'b1001101: c <= 9'b100100001;
				8'b111111: c <= 9'b10101100;
				8'b1101110: c <= 9'b111100111;
				8'b1111011: c <= 9'b11010101;
				8'b1001011: c <= 9'b101101001;
				8'b1101111: c <= 9'b1010001;
				8'b1101000: c <= 9'b1000010;
				8'b101100: c <= 9'b111110011;
				8'b100100: c <= 9'b100000111;
				8'b1111000: c <= 9'b111111;
				8'b1000101: c <= 9'b100110101;
				8'b1011001: c <= 9'b101011010;
				8'b110100: c <= 9'b101110111;
				8'b1111001: c <= 9'b110001;
				8'b1110001: c <= 9'b1010000;
				8'b1001111: c <= 9'b11111101;
				8'b1100101: c <= 9'b11100001;
				8'b1111110: c <= 9'b1010111;
				8'b1111100: c <= 9'b101001011;
				8'b1010110: c <= 9'b11011100;
				8'b110010: c <= 9'b101010000;
				8'b1101101: c <= 9'b11100000;
				8'b100011: c <= 9'b111011011;
				8'b1110101: c <= 9'b1110011;
				8'b1111101: c <= 9'b100110101;
				8'b101001: c <= 9'b100100101;
				8'b1010010: c <= 9'b111100011;
				8'b1011000: c <= 9'b101100;
				8'b101110: c <= 9'b111100100;
				8'b1000001: c <= 9'b11001110;
				default: c <= 9'b0;
			endcase
			9'b100011100 : case(di)
				8'b1000011: c <= 9'b10110;
				8'b101000: c <= 9'b1000;
				8'b111010: c <= 9'b101;
				8'b110110: c <= 9'b100110101;
				8'b1100100: c <= 9'b100000001;
				8'b1000000: c <= 9'b111000110;
				8'b1110110: c <= 9'b1101101;
				8'b100101: c <= 9'b10001010;
				8'b101111: c <= 9'b111000000;
				8'b100110: c <= 9'b1010101;
				8'b1100011: c <= 9'b1101001;
				8'b1001000: c <= 9'b10000110;
				8'b111000: c <= 9'b11000;
				8'b110001: c <= 9'b100010111;
				8'b1010111: c <= 9'b10111000;
				8'b1001110: c <= 9'b100110110;
				8'b1101010: c <= 9'b10000001;
				8'b1001001: c <= 9'b11011101;
				8'b1100000: c <= 9'b1011;
				8'b110111: c <= 9'b101110010;
				8'b1011101: c <= 9'b10010011;
				8'b1011011: c <= 9'b11000111;
				8'b111001: c <= 9'b11110001;
				8'b1001010: c <= 9'b10001100;
				8'b110011: c <= 9'b10010;
				8'b1101100: c <= 9'b110001100;
				8'b1110111: c <= 9'b100000010;
				8'b101011: c <= 9'b111100001;
				8'b1101011: c <= 9'b11001110;
				8'b111100: c <= 9'b11110100;
				8'b1000111: c <= 9'b1101010;
				8'b1011111: c <= 9'b100100001;
				8'b1110100: c <= 9'b110100110;
				8'b101101: c <= 9'b11101001;
				8'b1010011: c <= 9'b111101101;
				8'b1100001: c <= 9'b10011111;
				8'b110101: c <= 9'b110011010;
				8'b1000100: c <= 9'b11110110;
				8'b1010001: c <= 9'b110010111;
				8'b1010100: c <= 9'b1100010;
				8'b1100110: c <= 9'b100011010;
				8'b101010: c <= 9'b10010;
				8'b1011110: c <= 9'b100100111;
				8'b1100111: c <= 9'b1110101;
				8'b1011010: c <= 9'b11001110;
				8'b1000010: c <= 9'b100101111;
				8'b111101: c <= 9'b10100011;
				8'b110000: c <= 9'b100001010;
				8'b111110: c <= 9'b10001001;
				8'b1100010: c <= 9'b10101;
				8'b1110000: c <= 9'b110000110;
				8'b1101001: c <= 9'b110111010;
				8'b1110011: c <= 9'b110100;
				8'b1001100: c <= 9'b110100100;
				8'b100001: c <= 9'b11110;
				8'b1000110: c <= 9'b111101111;
				8'b1110010: c <= 9'b11010010;
				8'b1010000: c <= 9'b110111010;
				8'b1111010: c <= 9'b100001100;
				8'b1010101: c <= 9'b101100110;
				8'b111011: c <= 9'b10011000;
				8'b1001101: c <= 9'b10001000;
				8'b111111: c <= 9'b110100110;
				8'b1101110: c <= 9'b101101111;
				8'b1111011: c <= 9'b111011100;
				8'b1001011: c <= 9'b101110011;
				8'b1101111: c <= 9'b111001;
				8'b1101000: c <= 9'b110000101;
				8'b101100: c <= 9'b101011111;
				8'b100100: c <= 9'b11110001;
				8'b1111000: c <= 9'b1111010;
				8'b1000101: c <= 9'b10000011;
				8'b1011001: c <= 9'b110101101;
				8'b110100: c <= 9'b1110111;
				8'b1111001: c <= 9'b1011011;
				8'b1110001: c <= 9'b111001100;
				8'b1001111: c <= 9'b11001111;
				8'b1100101: c <= 9'b101000010;
				8'b1111110: c <= 9'b11000011;
				8'b1111100: c <= 9'b100101000;
				8'b1010110: c <= 9'b1101101;
				8'b110010: c <= 9'b11110100;
				8'b1101101: c <= 9'b10110;
				8'b100011: c <= 9'b101010100;
				8'b1110101: c <= 9'b10111000;
				8'b1111101: c <= 9'b100101010;
				8'b101001: c <= 9'b1100000;
				8'b1010010: c <= 9'b110100001;
				8'b1011000: c <= 9'b11010111;
				8'b101110: c <= 9'b100011000;
				8'b1000001: c <= 9'b110001110;
				default: c <= 9'b0;
			endcase
			9'b101011110 : case(di)
				8'b1000011: c <= 9'b100001011;
				8'b101000: c <= 9'b11100110;
				8'b111010: c <= 9'b1100100;
				8'b110110: c <= 9'b100011111;
				8'b1100100: c <= 9'b101011011;
				8'b1000000: c <= 9'b100111000;
				8'b1110110: c <= 9'b100010101;
				8'b100101: c <= 9'b1001111;
				8'b101111: c <= 9'b10101000;
				8'b100110: c <= 9'b1101000;
				8'b1100011: c <= 9'b11011;
				8'b1001000: c <= 9'b10011000;
				8'b111000: c <= 9'b111111010;
				8'b110001: c <= 9'b100001001;
				8'b1010111: c <= 9'b111101111;
				8'b1001110: c <= 9'b101100101;
				8'b1101010: c <= 9'b11011011;
				8'b1001001: c <= 9'b1100;
				8'b1100000: c <= 9'b110001001;
				8'b110111: c <= 9'b101010100;
				8'b1011101: c <= 9'b11100111;
				8'b1011011: c <= 9'b1010110;
				8'b111001: c <= 9'b111000;
				8'b1001010: c <= 9'b11010101;
				8'b110011: c <= 9'b1010101;
				8'b1101100: c <= 9'b11111011;
				8'b1110111: c <= 9'b100111001;
				8'b101011: c <= 9'b100110000;
				8'b1101011: c <= 9'b110100101;
				8'b111100: c <= 9'b1010010;
				8'b1000111: c <= 9'b100101010;
				8'b1011111: c <= 9'b100010000;
				8'b1110100: c <= 9'b11100101;
				8'b101101: c <= 9'b100110000;
				8'b1010011: c <= 9'b111011100;
				8'b1100001: c <= 9'b100000000;
				8'b110101: c <= 9'b101010;
				8'b1000100: c <= 9'b101;
				8'b1010001: c <= 9'b1110100;
				8'b1010100: c <= 9'b101010011;
				8'b1100110: c <= 9'b11111100;
				8'b101010: c <= 9'b1001111;
				8'b1011110: c <= 9'b111111101;
				8'b1100111: c <= 9'b110100100;
				8'b1011010: c <= 9'b110000101;
				8'b1000010: c <= 9'b11110001;
				8'b111101: c <= 9'b101110001;
				8'b110000: c <= 9'b11110101;
				8'b111110: c <= 9'b10010101;
				8'b1100010: c <= 9'b100100;
				8'b1110000: c <= 9'b10010110;
				8'b1101001: c <= 9'b1110001;
				8'b1110011: c <= 9'b10010110;
				8'b1001100: c <= 9'b1100011;
				8'b100001: c <= 9'b11110110;
				8'b1000110: c <= 9'b111101001;
				8'b1110010: c <= 9'b110001001;
				8'b1010000: c <= 9'b1110001;
				8'b1111010: c <= 9'b1011001;
				8'b1010101: c <= 9'b10000111;
				8'b111011: c <= 9'b110101;
				8'b1001101: c <= 9'b11100;
				8'b111111: c <= 9'b11000100;
				8'b1101110: c <= 9'b101001010;
				8'b1111011: c <= 9'b11101011;
				8'b1001011: c <= 9'b11111011;
				8'b1101111: c <= 9'b110101001;
				8'b1101000: c <= 9'b11110001;
				8'b101100: c <= 9'b101110001;
				8'b100100: c <= 9'b1011100;
				8'b1111000: c <= 9'b110001000;
				8'b1000101: c <= 9'b1110001;
				8'b1011001: c <= 9'b1011001;
				8'b110100: c <= 9'b111000100;
				8'b1111001: c <= 9'b10010110;
				8'b1110001: c <= 9'b110100000;
				8'b1001111: c <= 9'b11111000;
				8'b1100101: c <= 9'b10000;
				8'b1111110: c <= 9'b110011110;
				8'b1111100: c <= 9'b1000010;
				8'b1010110: c <= 9'b10011100;
				8'b110010: c <= 9'b11001111;
				8'b1101101: c <= 9'b11111011;
				8'b100011: c <= 9'b111000101;
				8'b1110101: c <= 9'b101101000;
				8'b1111101: c <= 9'b10000000;
				8'b101001: c <= 9'b110110100;
				8'b1010010: c <= 9'b10001000;
				8'b1011000: c <= 9'b110011010;
				8'b101110: c <= 9'b101100001;
				8'b1000001: c <= 9'b101100111;
				default: c <= 9'b0;
			endcase
			9'b11001101 : case(di)
				8'b1000011: c <= 9'b110000010;
				8'b101000: c <= 9'b1001101;
				8'b111010: c <= 9'b111111011;
				8'b110110: c <= 9'b11000000;
				8'b1100100: c <= 9'b111010;
				8'b1000000: c <= 9'b11100111;
				8'b1110110: c <= 9'b100101100;
				8'b100101: c <= 9'b10101000;
				8'b101111: c <= 9'b101101;
				8'b100110: c <= 9'b100110000;
				8'b1100011: c <= 9'b111111101;
				8'b1001000: c <= 9'b100101;
				8'b111000: c <= 9'b101110110;
				8'b110001: c <= 9'b101010001;
				8'b1010111: c <= 9'b10010;
				8'b1001110: c <= 9'b101111000;
				8'b1101010: c <= 9'b100100101;
				8'b1001001: c <= 9'b101011010;
				8'b1100000: c <= 9'b1011;
				8'b110111: c <= 9'b111101001;
				8'b1011101: c <= 9'b100111110;
				8'b1011011: c <= 9'b10010000;
				8'b111001: c <= 9'b110111111;
				8'b1001010: c <= 9'b110111;
				8'b110011: c <= 9'b10000111;
				8'b1101100: c <= 9'b100010110;
				8'b1110111: c <= 9'b1011011;
				8'b101011: c <= 9'b100010011;
				8'b1101011: c <= 9'b10101;
				8'b111100: c <= 9'b100001110;
				8'b1000111: c <= 9'b110001010;
				8'b1011111: c <= 9'b100100111;
				8'b1110100: c <= 9'b10000101;
				8'b101101: c <= 9'b110001101;
				8'b1010011: c <= 9'b10101;
				8'b1100001: c <= 9'b111110101;
				8'b110101: c <= 9'b11001010;
				8'b1000100: c <= 9'b110011010;
				8'b1010001: c <= 9'b111;
				8'b1010100: c <= 9'b11100100;
				8'b1100110: c <= 9'b10100000;
				8'b101010: c <= 9'b110110100;
				8'b1011110: c <= 9'b110110010;
				8'b1100111: c <= 9'b100100;
				8'b1011010: c <= 9'b1110;
				8'b1000010: c <= 9'b111100;
				8'b111101: c <= 9'b11011010;
				8'b110000: c <= 9'b100001110;
				8'b111110: c <= 9'b101001010;
				8'b1100010: c <= 9'b100011000;
				8'b1110000: c <= 9'b101000101;
				8'b1101001: c <= 9'b100010010;
				8'b1110011: c <= 9'b111000110;
				8'b1001100: c <= 9'b10110;
				8'b100001: c <= 9'b11111010;
				8'b1000110: c <= 9'b111111001;
				8'b1110010: c <= 9'b101011010;
				8'b1010000: c <= 9'b100111001;
				8'b1111010: c <= 9'b110000111;
				8'b1010101: c <= 9'b10111111;
				8'b111011: c <= 9'b101010101;
				8'b1001101: c <= 9'b110100010;
				8'b111111: c <= 9'b11011;
				8'b1101110: c <= 9'b1100011;
				8'b1111011: c <= 9'b111100;
				8'b1001011: c <= 9'b111011111;
				8'b1101111: c <= 9'b1010000;
				8'b1101000: c <= 9'b101001011;
				8'b101100: c <= 9'b1111010;
				8'b100100: c <= 9'b1;
				8'b1111000: c <= 9'b10011010;
				8'b1000101: c <= 9'b1110111;
				8'b1011001: c <= 9'b11100111;
				8'b110100: c <= 9'b110010001;
				8'b1111001: c <= 9'b101011;
				8'b1110001: c <= 9'b111111000;
				8'b1001111: c <= 9'b100110100;
				8'b1100101: c <= 9'b11111100;
				8'b1111110: c <= 9'b1110001;
				8'b1111100: c <= 9'b100110100;
				8'b1010110: c <= 9'b110110100;
				8'b110010: c <= 9'b100100110;
				8'b1101101: c <= 9'b11001010;
				8'b100011: c <= 9'b11111010;
				8'b1110101: c <= 9'b111100100;
				8'b1111101: c <= 9'b10010101;
				8'b101001: c <= 9'b1010110;
				8'b1010010: c <= 9'b1001101;
				8'b1011000: c <= 9'b11010111;
				8'b101110: c <= 9'b1000110;
				8'b1000001: c <= 9'b1111111;
				default: c <= 9'b0;
			endcase
			9'b10100011 : case(di)
				8'b1000011: c <= 9'b101100010;
				8'b101000: c <= 9'b10001000;
				8'b111010: c <= 9'b110100111;
				8'b110110: c <= 9'b101001100;
				8'b1100100: c <= 9'b110010101;
				8'b1000000: c <= 9'b11110100;
				8'b1110110: c <= 9'b11000;
				8'b100101: c <= 9'b100101100;
				8'b101111: c <= 9'b110001111;
				8'b100110: c <= 9'b100010;
				8'b1100011: c <= 9'b101010111;
				8'b1001000: c <= 9'b100000100;
				8'b111000: c <= 9'b1110101;
				8'b110001: c <= 9'b110100101;
				8'b1010111: c <= 9'b101111001;
				8'b1001110: c <= 9'b11000010;
				8'b1101010: c <= 9'b11011100;
				8'b1001001: c <= 9'b11010100;
				8'b1100000: c <= 9'b10001001;
				8'b110111: c <= 9'b1111010;
				8'b1011101: c <= 9'b11000;
				8'b1011011: c <= 9'b101000111;
				8'b111001: c <= 9'b1010011;
				8'b1001010: c <= 9'b1011000;
				8'b110011: c <= 9'b111100;
				8'b1101100: c <= 9'b1011100;
				8'b1110111: c <= 9'b110011100;
				8'b101011: c <= 9'b100001110;
				8'b1101011: c <= 9'b1011100;
				8'b111100: c <= 9'b111100111;
				8'b1000111: c <= 9'b111011110;
				8'b1011111: c <= 9'b1000110;
				8'b1110100: c <= 9'b100010000;
				8'b101101: c <= 9'b110010011;
				8'b1010011: c <= 9'b111011010;
				8'b1100001: c <= 9'b110101111;
				8'b110101: c <= 9'b100111010;
				8'b1000100: c <= 9'b111101110;
				8'b1010001: c <= 9'b101110001;
				8'b1010100: c <= 9'b101100;
				8'b1100110: c <= 9'b1010010;
				8'b101010: c <= 9'b111000;
				8'b1011110: c <= 9'b100101011;
				8'b1100111: c <= 9'b11100111;
				8'b1011010: c <= 9'b1001001;
				8'b1000010: c <= 9'b110011111;
				8'b111101: c <= 9'b1001;
				8'b110000: c <= 9'b110100011;
				8'b111110: c <= 9'b100111011;
				8'b1100010: c <= 9'b10010100;
				8'b1110000: c <= 9'b100001001;
				8'b1101001: c <= 9'b10101110;
				8'b1110011: c <= 9'b100111010;
				8'b1001100: c <= 9'b101001100;
				8'b100001: c <= 9'b100111111;
				8'b1000110: c <= 9'b101110000;
				8'b1110010: c <= 9'b100111001;
				8'b1010000: c <= 9'b111000100;
				8'b1111010: c <= 9'b10111111;
				8'b1010101: c <= 9'b10000;
				8'b111011: c <= 9'b101010101;
				8'b1001101: c <= 9'b101010000;
				8'b111111: c <= 9'b100011001;
				8'b1101110: c <= 9'b110101100;
				8'b1111011: c <= 9'b101000001;
				8'b1001011: c <= 9'b101011010;
				8'b1101111: c <= 9'b10010000;
				8'b1101000: c <= 9'b100001101;
				8'b101100: c <= 9'b11100001;
				8'b100100: c <= 9'b11001011;
				8'b1111000: c <= 9'b110101111;
				8'b1000101: c <= 9'b111011011;
				8'b1011001: c <= 9'b1000110;
				8'b110100: c <= 9'b100011000;
				8'b1111001: c <= 9'b10000010;
				8'b1110001: c <= 9'b11000011;
				8'b1001111: c <= 9'b100110000;
				8'b1100101: c <= 9'b100011011;
				8'b1111110: c <= 9'b10001111;
				8'b1111100: c <= 9'b11001001;
				8'b1010110: c <= 9'b110110;
				8'b110010: c <= 9'b11011010;
				8'b1101101: c <= 9'b101100101;
				8'b100011: c <= 9'b111110000;
				8'b1110101: c <= 9'b10110;
				8'b1111101: c <= 9'b11110;
				8'b101001: c <= 9'b100000001;
				8'b1010010: c <= 9'b101101;
				8'b1011000: c <= 9'b101101001;
				8'b101110: c <= 9'b10101101;
				8'b1000001: c <= 9'b100001111;
				default: c <= 9'b0;
			endcase
			9'b101110000 : case(di)
				8'b1000011: c <= 9'b11000011;
				8'b101000: c <= 9'b10111000;
				8'b111010: c <= 9'b101101000;
				8'b110110: c <= 9'b100001011;
				8'b1100100: c <= 9'b1110111;
				8'b1000000: c <= 9'b101101101;
				8'b1110110: c <= 9'b1010101;
				8'b100101: c <= 9'b100010111;
				8'b101111: c <= 9'b101110110;
				8'b100110: c <= 9'b1010110;
				8'b1100011: c <= 9'b11111101;
				8'b1001000: c <= 9'b111101;
				8'b111000: c <= 9'b110111001;
				8'b110001: c <= 9'b100110010;
				8'b1010111: c <= 9'b111100111;
				8'b1001110: c <= 9'b100011000;
				8'b1101010: c <= 9'b1100111;
				8'b1001001: c <= 9'b11101111;
				8'b1100000: c <= 9'b1000110;
				8'b110111: c <= 9'b111100000;
				8'b1011101: c <= 9'b100101001;
				8'b1011011: c <= 9'b111010100;
				8'b111001: c <= 9'b10110010;
				8'b1001010: c <= 9'b100111011;
				8'b110011: c <= 9'b100000101;
				8'b1101100: c <= 9'b110101111;
				8'b1110111: c <= 9'b1001101;
				8'b101011: c <= 9'b1001110;
				8'b1101011: c <= 9'b10000010;
				8'b111100: c <= 9'b10100101;
				8'b1000111: c <= 9'b11110011;
				8'b1011111: c <= 9'b110010010;
				8'b1110100: c <= 9'b111001010;
				8'b101101: c <= 9'b11100001;
				8'b1010011: c <= 9'b100100;
				8'b1100001: c <= 9'b10100100;
				8'b110101: c <= 9'b111000110;
				8'b1000100: c <= 9'b11101001;
				8'b1010001: c <= 9'b101010000;
				8'b1010100: c <= 9'b110011101;
				8'b1100110: c <= 9'b110101011;
				8'b101010: c <= 9'b110011;
				8'b1011110: c <= 9'b110110100;
				8'b1100111: c <= 9'b101000110;
				8'b1011010: c <= 9'b101010010;
				8'b1000010: c <= 9'b100010110;
				8'b111101: c <= 9'b11000011;
				8'b110000: c <= 9'b110110010;
				8'b111110: c <= 9'b100001010;
				8'b1100010: c <= 9'b1000010;
				8'b1110000: c <= 9'b100001;
				8'b1101001: c <= 9'b110100110;
				8'b1110011: c <= 9'b101010000;
				8'b1001100: c <= 9'b1111100;
				8'b100001: c <= 9'b101101011;
				8'b1000110: c <= 9'b100000101;
				8'b1110010: c <= 9'b11110011;
				8'b1010000: c <= 9'b10010100;
				8'b1111010: c <= 9'b11101111;
				8'b1010101: c <= 9'b101010;
				8'b111011: c <= 9'b111000;
				8'b1001101: c <= 9'b100101101;
				8'b111111: c <= 9'b110101001;
				8'b1101110: c <= 9'b111100111;
				8'b1111011: c <= 9'b1101101;
				8'b1001011: c <= 9'b111001;
				8'b1101111: c <= 9'b101101110;
				8'b1101000: c <= 9'b11101;
				8'b101100: c <= 9'b10100010;
				8'b100100: c <= 9'b100111011;
				8'b1111000: c <= 9'b111100;
				8'b1000101: c <= 9'b1010010;
				8'b1011001: c <= 9'b100000100;
				8'b110100: c <= 9'b100011010;
				8'b1111001: c <= 9'b110;
				8'b1110001: c <= 9'b11011010;
				8'b1001111: c <= 9'b101100110;
				8'b1100101: c <= 9'b111011011;
				8'b1111110: c <= 9'b111011111;
				8'b1111100: c <= 9'b1001000;
				8'b1010110: c <= 9'b100001101;
				8'b110010: c <= 9'b100111000;
				8'b1101101: c <= 9'b100101111;
				8'b100011: c <= 9'b1001001;
				8'b1110101: c <= 9'b111000100;
				8'b1111101: c <= 9'b1011011;
				8'b101001: c <= 9'b100010110;
				8'b1010010: c <= 9'b101000010;
				8'b1011000: c <= 9'b111100010;
				8'b101110: c <= 9'b11100101;
				8'b1000001: c <= 9'b111010001;
				default: c <= 9'b0;
			endcase
			9'b111000010 : case(di)
				8'b1000011: c <= 9'b111000100;
				8'b101000: c <= 9'b10101100;
				8'b111010: c <= 9'b100010110;
				8'b110110: c <= 9'b11100110;
				8'b1100100: c <= 9'b10101010;
				8'b1000000: c <= 9'b111010110;
				8'b1110110: c <= 9'b100;
				8'b100101: c <= 9'b11011101;
				8'b101111: c <= 9'b110000101;
				8'b100110: c <= 9'b1000111;
				8'b1100011: c <= 9'b100001110;
				8'b1001000: c <= 9'b100011000;
				8'b111000: c <= 9'b10011001;
				8'b110001: c <= 9'b100;
				8'b1010111: c <= 9'b110;
				8'b1001110: c <= 9'b10110001;
				8'b1101010: c <= 9'b1100101;
				8'b1001001: c <= 9'b110011111;
				8'b1100000: c <= 9'b10100110;
				8'b110111: c <= 9'b110111;
				8'b1011101: c <= 9'b1111100;
				8'b1011011: c <= 9'b110000101;
				8'b111001: c <= 9'b110010;
				8'b1001010: c <= 9'b111111110;
				8'b110011: c <= 9'b111000011;
				8'b1101100: c <= 9'b101010000;
				8'b1110111: c <= 9'b100101111;
				8'b101011: c <= 9'b10000000;
				8'b1101011: c <= 9'b101111010;
				8'b111100: c <= 9'b101010000;
				8'b1000111: c <= 9'b111001010;
				8'b1011111: c <= 9'b100011000;
				8'b1110100: c <= 9'b101111001;
				8'b101101: c <= 9'b10000001;
				8'b1010011: c <= 9'b111101110;
				8'b1100001: c <= 9'b100111101;
				8'b110101: c <= 9'b11011101;
				8'b1000100: c <= 9'b100101000;
				8'b1010001: c <= 9'b111100110;
				8'b1010100: c <= 9'b110101100;
				8'b1100110: c <= 9'b100111111;
				8'b101010: c <= 9'b110011;
				8'b1011110: c <= 9'b100101110;
				8'b1100111: c <= 9'b10110010;
				8'b1011010: c <= 9'b1110100;
				8'b1000010: c <= 9'b100100000;
				8'b111101: c <= 9'b11001101;
				8'b110000: c <= 9'b111001001;
				8'b111110: c <= 9'b110011111;
				8'b1100010: c <= 9'b10001110;
				8'b1110000: c <= 9'b11101000;
				8'b1101001: c <= 9'b111010010;
				8'b1110011: c <= 9'b10010100;
				8'b1001100: c <= 9'b101101001;
				8'b100001: c <= 9'b11110010;
				8'b1000110: c <= 9'b10100111;
				8'b1110010: c <= 9'b101011000;
				8'b1010000: c <= 9'b1010001;
				8'b1111010: c <= 9'b110101110;
				8'b1010101: c <= 9'b110010101;
				8'b111011: c <= 9'b101000101;
				8'b1001101: c <= 9'b100001011;
				8'b111111: c <= 9'b100110100;
				8'b1101110: c <= 9'b1011110;
				8'b1111011: c <= 9'b101011010;
				8'b1001011: c <= 9'b111001100;
				8'b1101111: c <= 9'b100001;
				8'b1101000: c <= 9'b100010011;
				8'b101100: c <= 9'b10011000;
				8'b100100: c <= 9'b111000110;
				8'b1111000: c <= 9'b101000111;
				8'b1000101: c <= 9'b1000111;
				8'b1011001: c <= 9'b110111;
				8'b110100: c <= 9'b110110011;
				8'b1111001: c <= 9'b111010001;
				8'b1110001: c <= 9'b111100010;
				8'b1001111: c <= 9'b10010101;
				8'b1100101: c <= 9'b111111011;
				8'b1111110: c <= 9'b1001;
				8'b1111100: c <= 9'b101111000;
				8'b1010110: c <= 9'b11001111;
				8'b110010: c <= 9'b101010;
				8'b1101101: c <= 9'b110000110;
				8'b100011: c <= 9'b111001111;
				8'b1110101: c <= 9'b10111100;
				8'b1111101: c <= 9'b10111000;
				8'b101001: c <= 9'b110110011;
				8'b1010010: c <= 9'b1011001;
				8'b1011000: c <= 9'b100001101;
				8'b101110: c <= 9'b110011011;
				8'b1000001: c <= 9'b100111101;
				default: c <= 9'b0;
			endcase
			9'b101101111 : case(di)
				8'b1000011: c <= 9'b101001000;
				8'b101000: c <= 9'b1111110;
				8'b111010: c <= 9'b110110010;
				8'b110110: c <= 9'b11101;
				8'b1100100: c <= 9'b101010;
				8'b1000000: c <= 9'b10111111;
				8'b1110110: c <= 9'b10110101;
				8'b100101: c <= 9'b11000100;
				8'b101111: c <= 9'b10111;
				8'b100110: c <= 9'b101000010;
				8'b1100011: c <= 9'b101101101;
				8'b1001000: c <= 9'b1100;
				8'b111000: c <= 9'b100001;
				8'b110001: c <= 9'b101100010;
				8'b1010111: c <= 9'b110100000;
				8'b1001110: c <= 9'b111101100;
				8'b1101010: c <= 9'b10011000;
				8'b1001001: c <= 9'b11010000;
				8'b1100000: c <= 9'b110101;
				8'b110111: c <= 9'b11100001;
				8'b1011101: c <= 9'b100110100;
				8'b1011011: c <= 9'b1011;
				8'b111001: c <= 9'b100;
				8'b1001010: c <= 9'b10110011;
				8'b110011: c <= 9'b110011001;
				8'b1101100: c <= 9'b10111001;
				8'b1110111: c <= 9'b110110111;
				8'b101011: c <= 9'b11001;
				8'b1101011: c <= 9'b111;
				8'b111100: c <= 9'b100010;
				8'b1000111: c <= 9'b11010011;
				8'b1011111: c <= 9'b11010100;
				8'b1110100: c <= 9'b1000010;
				8'b101101: c <= 9'b11101000;
				8'b1010011: c <= 9'b10000111;
				8'b1100001: c <= 9'b10100110;
				8'b110101: c <= 9'b100011;
				8'b1000100: c <= 9'b101111010;
				8'b1010001: c <= 9'b1011001;
				8'b1010100: c <= 9'b111000000;
				8'b1100110: c <= 9'b10011101;
				8'b101010: c <= 9'b10001111;
				8'b1011110: c <= 9'b111111;
				8'b1100111: c <= 9'b111011111;
				8'b1011010: c <= 9'b1010110;
				8'b1000010: c <= 9'b110101010;
				8'b111101: c <= 9'b11011;
				8'b110000: c <= 9'b1101010;
				8'b111110: c <= 9'b111001101;
				8'b1100010: c <= 9'b100001100;
				8'b1110000: c <= 9'b100010100;
				8'b1101001: c <= 9'b111011010;
				8'b1110011: c <= 9'b101000100;
				8'b1001100: c <= 9'b100011010;
				8'b100001: c <= 9'b101010;
				8'b1000110: c <= 9'b11000000;
				8'b1110010: c <= 9'b11001001;
				8'b1010000: c <= 9'b111;
				8'b1111010: c <= 9'b110;
				8'b1010101: c <= 9'b110100010;
				8'b111011: c <= 9'b101000010;
				8'b1001101: c <= 9'b1100011;
				8'b111111: c <= 9'b11010010;
				8'b1101110: c <= 9'b11010101;
				8'b1111011: c <= 9'b1101110;
				8'b1001011: c <= 9'b100011;
				8'b1101111: c <= 9'b111001111;
				8'b1101000: c <= 9'b10011001;
				8'b101100: c <= 9'b100011101;
				8'b100100: c <= 9'b1100000;
				8'b1111000: c <= 9'b11110100;
				8'b1000101: c <= 9'b100011100;
				8'b1011001: c <= 9'b11011;
				8'b110100: c <= 9'b100100011;
				8'b1111001: c <= 9'b111111110;
				8'b1110001: c <= 9'b101101;
				8'b1001111: c <= 9'b111100010;
				8'b1100101: c <= 9'b101010011;
				8'b1111110: c <= 9'b110001101;
				8'b1111100: c <= 9'b10100101;
				8'b1010110: c <= 9'b101010110;
				8'b110010: c <= 9'b111100111;
				8'b1101101: c <= 9'b10010100;
				8'b100011: c <= 9'b100;
				8'b1110101: c <= 9'b111001001;
				8'b1111101: c <= 9'b10010000;
				8'b101001: c <= 9'b10100011;
				8'b1010010: c <= 9'b11100;
				8'b1011000: c <= 9'b100101010;
				8'b101110: c <= 9'b100001010;
				8'b1000001: c <= 9'b110101111;
				default: c <= 9'b0;
			endcase
			9'b10011010 : case(di)
				8'b1000011: c <= 9'b1001110;
				8'b101000: c <= 9'b11001000;
				8'b111010: c <= 9'b101110110;
				8'b110110: c <= 9'b10011100;
				8'b1100100: c <= 9'b100010001;
				8'b1000000: c <= 9'b1001100;
				8'b1110110: c <= 9'b11000011;
				8'b100101: c <= 9'b111011111;
				8'b101111: c <= 9'b111011011;
				8'b100110: c <= 9'b101101001;
				8'b1100011: c <= 9'b10011100;
				8'b1001000: c <= 9'b10000110;
				8'b111000: c <= 9'b110000;
				8'b110001: c <= 9'b100101011;
				8'b1010111: c <= 9'b100010001;
				8'b1001110: c <= 9'b10110;
				8'b1101010: c <= 9'b101000;
				8'b1001001: c <= 9'b1001100;
				8'b1100000: c <= 9'b110010110;
				8'b110111: c <= 9'b101000111;
				8'b1011101: c <= 9'b10001000;
				8'b1011011: c <= 9'b11100;
				8'b111001: c <= 9'b1110;
				8'b1001010: c <= 9'b111100000;
				8'b110011: c <= 9'b101000100;
				8'b1101100: c <= 9'b11000100;
				8'b1110111: c <= 9'b101101111;
				8'b101011: c <= 9'b101000010;
				8'b1101011: c <= 9'b110010111;
				8'b111100: c <= 9'b111001100;
				8'b1000111: c <= 9'b101001011;
				8'b1011111: c <= 9'b11001100;
				8'b1110100: c <= 9'b110000;
				8'b101101: c <= 9'b11010000;
				8'b1010011: c <= 9'b101101001;
				8'b1100001: c <= 9'b110111011;
				8'b110101: c <= 9'b10011;
				8'b1000100: c <= 9'b11111110;
				8'b1010001: c <= 9'b101001011;
				8'b1010100: c <= 9'b100000100;
				8'b1100110: c <= 9'b1000011;
				8'b101010: c <= 9'b100110000;
				8'b1011110: c <= 9'b1100010;
				8'b1100111: c <= 9'b11001001;
				8'b1011010: c <= 9'b111000110;
				8'b1000010: c <= 9'b1111001;
				8'b111101: c <= 9'b111001011;
				8'b110000: c <= 9'b111011100;
				8'b111110: c <= 9'b10111111;
				8'b1100010: c <= 9'b110111000;
				8'b1110000: c <= 9'b11010;
				8'b1101001: c <= 9'b11010011;
				8'b1110011: c <= 9'b1001;
				8'b1001100: c <= 9'b10101000;
				8'b100001: c <= 9'b101001011;
				8'b1000110: c <= 9'b1101101;
				8'b1110010: c <= 9'b111000010;
				8'b1010000: c <= 9'b101111110;
				8'b1111010: c <= 9'b1101000;
				8'b1010101: c <= 9'b100110100;
				8'b111011: c <= 9'b10000011;
				8'b1001101: c <= 9'b10110001;
				8'b111111: c <= 9'b1101110;
				8'b1101110: c <= 9'b100110110;
				8'b1111011: c <= 9'b101110100;
				8'b1001011: c <= 9'b110000001;
				8'b1101111: c <= 9'b11001100;
				8'b1101000: c <= 9'b10010110;
				8'b101100: c <= 9'b111010000;
				8'b100100: c <= 9'b110011000;
				8'b1111000: c <= 9'b1100;
				8'b1000101: c <= 9'b100101111;
				8'b1011001: c <= 9'b11100101;
				8'b110100: c <= 9'b111011;
				8'b1111001: c <= 9'b100000101;
				8'b1110001: c <= 9'b1110001;
				8'b1001111: c <= 9'b11100011;
				8'b1100101: c <= 9'b111100110;
				8'b1111110: c <= 9'b100010011;
				8'b1111100: c <= 9'b100100000;
				8'b1010110: c <= 9'b10101001;
				8'b110010: c <= 9'b101000100;
				8'b1101101: c <= 9'b111011010;
				8'b100011: c <= 9'b10000101;
				8'b1110101: c <= 9'b11000000;
				8'b1111101: c <= 9'b111011;
				8'b101001: c <= 9'b100010;
				8'b1010010: c <= 9'b101011111;
				8'b1011000: c <= 9'b1001010;
				8'b101110: c <= 9'b111100000;
				8'b1000001: c <= 9'b10010;
				default: c <= 9'b0;
			endcase
			9'b11001100 : case(di)
				8'b1000011: c <= 9'b11100000;
				8'b101000: c <= 9'b110101101;
				8'b111010: c <= 9'b101001010;
				8'b110110: c <= 9'b1100011;
				8'b1100100: c <= 9'b101011000;
				8'b1000000: c <= 9'b110101101;
				8'b1110110: c <= 9'b10101110;
				8'b100101: c <= 9'b10111010;
				8'b101111: c <= 9'b110100101;
				8'b100110: c <= 9'b1101010;
				8'b1100011: c <= 9'b1011;
				8'b1001000: c <= 9'b110;
				8'b111000: c <= 9'b101010100;
				8'b110001: c <= 9'b11010000;
				8'b1010111: c <= 9'b100101100;
				8'b1001110: c <= 9'b10010011;
				8'b1101010: c <= 9'b11110100;
				8'b1001001: c <= 9'b101010111;
				8'b1100000: c <= 9'b10;
				8'b110111: c <= 9'b111011101;
				8'b1011101: c <= 9'b111010111;
				8'b1011011: c <= 9'b111001;
				8'b111001: c <= 9'b101000010;
				8'b1001010: c <= 9'b10011111;
				8'b110011: c <= 9'b10100011;
				8'b1101100: c <= 9'b10011111;
				8'b1110111: c <= 9'b110001110;
				8'b101011: c <= 9'b110101011;
				8'b1101011: c <= 9'b101100111;
				8'b111100: c <= 9'b10111;
				8'b1000111: c <= 9'b111111011;
				8'b1011111: c <= 9'b100000100;
				8'b1110100: c <= 9'b110001;
				8'b101101: c <= 9'b100111111;
				8'b1010011: c <= 9'b10101100;
				8'b1100001: c <= 9'b10001011;
				8'b110101: c <= 9'b110101110;
				8'b1000100: c <= 9'b11100111;
				8'b1010001: c <= 9'b11110101;
				8'b1010100: c <= 9'b111011011;
				8'b1100110: c <= 9'b101001100;
				8'b101010: c <= 9'b11111110;
				8'b1011110: c <= 9'b100100111;
				8'b1100111: c <= 9'b11010;
				8'b1011010: c <= 9'b11000000;
				8'b1000010: c <= 9'b111001101;
				8'b111101: c <= 9'b1001111;
				8'b110000: c <= 9'b10010100;
				8'b111110: c <= 9'b110111;
				8'b1100010: c <= 9'b1100110;
				8'b1110000: c <= 9'b100111111;
				8'b1101001: c <= 9'b110011010;
				8'b1110011: c <= 9'b101100001;
				8'b1001100: c <= 9'b1110001;
				8'b100001: c <= 9'b111111001;
				8'b1000110: c <= 9'b11010;
				8'b1110010: c <= 9'b1011011;
				8'b1010000: c <= 9'b10111000;
				8'b1111010: c <= 9'b101000100;
				8'b1010101: c <= 9'b10111011;
				8'b111011: c <= 9'b100111001;
				8'b1001101: c <= 9'b110101110;
				8'b111111: c <= 9'b11010;
				8'b1101110: c <= 9'b100000010;
				8'b1111011: c <= 9'b111010010;
				8'b1001011: c <= 9'b101110110;
				8'b1101111: c <= 9'b110011011;
				8'b1101000: c <= 9'b1111011;
				8'b101100: c <= 9'b100100000;
				8'b100100: c <= 9'b10101111;
				8'b1111000: c <= 9'b111001000;
				8'b1000101: c <= 9'b101110000;
				8'b1011001: c <= 9'b10111110;
				8'b110100: c <= 9'b100001;
				8'b1111001: c <= 9'b101111010;
				8'b1110001: c <= 9'b111000100;
				8'b1001111: c <= 9'b101110000;
				8'b1100101: c <= 9'b11001101;
				8'b1111110: c <= 9'b100111001;
				8'b1111100: c <= 9'b1001001;
				8'b1010110: c <= 9'b110100001;
				8'b110010: c <= 9'b10111101;
				8'b1101101: c <= 9'b101010;
				8'b100011: c <= 9'b111010000;
				8'b1110101: c <= 9'b10101100;
				8'b1111101: c <= 9'b101000110;
				8'b101001: c <= 9'b10000011;
				8'b1010010: c <= 9'b10010001;
				8'b1011000: c <= 9'b110100110;
				8'b101110: c <= 9'b10010101;
				8'b1000001: c <= 9'b11011;
				default: c <= 9'b0;
			endcase
			9'b100100001 : case(di)
				8'b1000011: c <= 9'b111100010;
				8'b101000: c <= 9'b11000000;
				8'b111010: c <= 9'b1;
				8'b110110: c <= 9'b10000101;
				8'b1100100: c <= 9'b111011010;
				8'b1000000: c <= 9'b110010011;
				8'b1110110: c <= 9'b100100010;
				8'b100101: c <= 9'b101000010;
				8'b101111: c <= 9'b1111100;
				8'b100110: c <= 9'b100010000;
				8'b1100011: c <= 9'b11011010;
				8'b1001000: c <= 9'b100110111;
				8'b111000: c <= 9'b101111110;
				8'b110001: c <= 9'b101011011;
				8'b1010111: c <= 9'b11001111;
				8'b1001110: c <= 9'b10110100;
				8'b1101010: c <= 9'b110000011;
				8'b1001001: c <= 9'b10000110;
				8'b1100000: c <= 9'b10111110;
				8'b110111: c <= 9'b1010010;
				8'b1011101: c <= 9'b10001010;
				8'b1011011: c <= 9'b11111010;
				8'b111001: c <= 9'b10011010;
				8'b1001010: c <= 9'b110110111;
				8'b110011: c <= 9'b1001010;
				8'b1101100: c <= 9'b111011100;
				8'b1110111: c <= 9'b1001001;
				8'b101011: c <= 9'b100011011;
				8'b1101011: c <= 9'b10011100;
				8'b111100: c <= 9'b101010111;
				8'b1000111: c <= 9'b101101001;
				8'b1011111: c <= 9'b10110100;
				8'b1110100: c <= 9'b10101010;
				8'b101101: c <= 9'b101000010;
				8'b1010011: c <= 9'b10101000;
				8'b1100001: c <= 9'b101011011;
				8'b110101: c <= 9'b111100111;
				8'b1000100: c <= 9'b1000011;
				8'b1010001: c <= 9'b111100000;
				8'b1010100: c <= 9'b101010110;
				8'b1100110: c <= 9'b101010;
				8'b101010: c <= 9'b110011001;
				8'b1011110: c <= 9'b11110101;
				8'b1100111: c <= 9'b100000100;
				8'b1011010: c <= 9'b1101010;
				8'b1000010: c <= 9'b10101000;
				8'b111101: c <= 9'b10000101;
				8'b110000: c <= 9'b10100010;
				8'b111110: c <= 9'b110000110;
				8'b1100010: c <= 9'b11001111;
				8'b1110000: c <= 9'b11110100;
				8'b1101001: c <= 9'b100000111;
				8'b1110011: c <= 9'b110011100;
				8'b1001100: c <= 9'b110011010;
				8'b100001: c <= 9'b10010000;
				8'b1000110: c <= 9'b1000011;
				8'b1110010: c <= 9'b10001100;
				8'b1010000: c <= 9'b101110100;
				8'b1111010: c <= 9'b111010110;
				8'b1010101: c <= 9'b110101;
				8'b111011: c <= 9'b101001001;
				8'b1001101: c <= 9'b1111;
				8'b111111: c <= 9'b110001101;
				8'b1101110: c <= 9'b11110110;
				8'b1111011: c <= 9'b100101100;
				8'b1001011: c <= 9'b10011101;
				8'b1101111: c <= 9'b101001;
				8'b1101000: c <= 9'b10001101;
				8'b101100: c <= 9'b111011100;
				8'b100100: c <= 9'b1110001;
				8'b1111000: c <= 9'b101011000;
				8'b1000101: c <= 9'b100011111;
				8'b1011001: c <= 9'b110100;
				8'b110100: c <= 9'b1110100;
				8'b1111001: c <= 9'b100111010;
				8'b1110001: c <= 9'b111001100;
				8'b1001111: c <= 9'b100111001;
				8'b1100101: c <= 9'b1011111;
				8'b1111110: c <= 9'b100011101;
				8'b1111100: c <= 9'b1011011;
				8'b1010110: c <= 9'b1111111;
				8'b110010: c <= 9'b100100111;
				8'b1101101: c <= 9'b111111000;
				8'b100011: c <= 9'b10110110;
				8'b1110101: c <= 9'b110100011;
				8'b1111101: c <= 9'b1111100;
				8'b101001: c <= 9'b110111111;
				8'b1010010: c <= 9'b100100111;
				8'b1011000: c <= 9'b10100110;
				8'b101110: c <= 9'b111110110;
				8'b1000001: c <= 9'b11010011;
				default: c <= 9'b0;
			endcase
			9'b10010011 : case(di)
				8'b1000011: c <= 9'b111000100;
				8'b101000: c <= 9'b100101010;
				8'b111010: c <= 9'b11000010;
				8'b110110: c <= 9'b110001;
				8'b1100100: c <= 9'b101101010;
				8'b1000000: c <= 9'b110111;
				8'b1110110: c <= 9'b110010;
				8'b100101: c <= 9'b1101000;
				8'b101111: c <= 9'b111000100;
				8'b100110: c <= 9'b1111010;
				8'b1100011: c <= 9'b10010001;
				8'b1001000: c <= 9'b100101001;
				8'b111000: c <= 9'b1000010;
				8'b110001: c <= 9'b10010000;
				8'b1010111: c <= 9'b101110111;
				8'b1001110: c <= 9'b1110111;
				8'b1101010: c <= 9'b111000101;
				8'b1001001: c <= 9'b1010011;
				8'b1100000: c <= 9'b10001010;
				8'b110111: c <= 9'b100011010;
				8'b1011101: c <= 9'b110000001;
				8'b1011011: c <= 9'b101;
				8'b111001: c <= 9'b11101;
				8'b1001010: c <= 9'b111001111;
				8'b110011: c <= 9'b10011111;
				8'b1101100: c <= 9'b11011101;
				8'b1110111: c <= 9'b111011011;
				8'b101011: c <= 9'b111100100;
				8'b1101011: c <= 9'b100100000;
				8'b111100: c <= 9'b110010010;
				8'b1000111: c <= 9'b101101111;
				8'b1011111: c <= 9'b11010111;
				8'b1110100: c <= 9'b101110000;
				8'b101101: c <= 9'b1111100;
				8'b1010011: c <= 9'b1000101;
				8'b1100001: c <= 9'b101111111;
				8'b110101: c <= 9'b10000000;
				8'b1000100: c <= 9'b100011001;
				8'b1010001: c <= 9'b100100000;
				8'b1010100: c <= 9'b100101110;
				8'b1100110: c <= 9'b1011111;
				8'b101010: c <= 9'b1101;
				8'b1011110: c <= 9'b101111111;
				8'b1100111: c <= 9'b10011011;
				8'b1011010: c <= 9'b1110101;
				8'b1000010: c <= 9'b101011;
				8'b111101: c <= 9'b1110;
				8'b110000: c <= 9'b1100;
				8'b111110: c <= 9'b11110101;
				8'b1100010: c <= 9'b101110110;
				8'b1110000: c <= 9'b101110101;
				8'b1101001: c <= 9'b100100000;
				8'b1110011: c <= 9'b1001111;
				8'b1001100: c <= 9'b110100110;
				8'b100001: c <= 9'b110111011;
				8'b1000110: c <= 9'b11001011;
				8'b1110010: c <= 9'b111111001;
				8'b1010000: c <= 9'b111111111;
				8'b1111010: c <= 9'b11011001;
				8'b1010101: c <= 9'b10101101;
				8'b111011: c <= 9'b100001011;
				8'b1001101: c <= 9'b110100101;
				8'b111111: c <= 9'b1101;
				8'b1101110: c <= 9'b1110100;
				8'b1111011: c <= 9'b10000000;
				8'b1001011: c <= 9'b100010010;
				8'b1101111: c <= 9'b110111010;
				8'b1101000: c <= 9'b110110110;
				8'b101100: c <= 9'b10100000;
				8'b100100: c <= 9'b111111010;
				8'b1111000: c <= 9'b10100101;
				8'b1000101: c <= 9'b111111001;
				8'b1011001: c <= 9'b1000;
				8'b110100: c <= 9'b110100011;
				8'b1111001: c <= 9'b11010001;
				8'b1110001: c <= 9'b110101101;
				8'b1001111: c <= 9'b111000000;
				8'b1100101: c <= 9'b10000000;
				8'b1111110: c <= 9'b101000111;
				8'b1111100: c <= 9'b110011100;
				8'b1010110: c <= 9'b100111;
				8'b110010: c <= 9'b111000010;
				8'b1101101: c <= 9'b101001010;
				8'b100011: c <= 9'b101000;
				8'b1110101: c <= 9'b11010111;
				8'b1111101: c <= 9'b11001011;
				8'b101001: c <= 9'b111101;
				8'b1010010: c <= 9'b100000110;
				8'b1011000: c <= 9'b110001;
				8'b101110: c <= 9'b1101110;
				8'b1000001: c <= 9'b101111110;
				default: c <= 9'b0;
			endcase
			9'b111010000 : case(di)
				8'b1000011: c <= 9'b101111001;
				8'b101000: c <= 9'b110010;
				8'b111010: c <= 9'b101001100;
				8'b110110: c <= 9'b100100011;
				8'b1100100: c <= 9'b100000010;
				8'b1000000: c <= 9'b11110000;
				8'b1110110: c <= 9'b111011101;
				8'b100101: c <= 9'b10100101;
				8'b101111: c <= 9'b101010;
				8'b100110: c <= 9'b111111001;
				8'b1100011: c <= 9'b1000001;
				8'b1001000: c <= 9'b10001011;
				8'b111000: c <= 9'b100111101;
				8'b110001: c <= 9'b100011001;
				8'b1010111: c <= 9'b1010010;
				8'b1001110: c <= 9'b101000100;
				8'b1101010: c <= 9'b110011101;
				8'b1001001: c <= 9'b11000000;
				8'b1100000: c <= 9'b101111111;
				8'b110111: c <= 9'b100001001;
				8'b1011101: c <= 9'b101011001;
				8'b1011011: c <= 9'b11010010;
				8'b111001: c <= 9'b100101101;
				8'b1001010: c <= 9'b100011111;
				8'b110011: c <= 9'b111001111;
				8'b1101100: c <= 9'b11000;
				8'b1110111: c <= 9'b100011001;
				8'b101011: c <= 9'b100100;
				8'b1101011: c <= 9'b10101;
				8'b111100: c <= 9'b10010001;
				8'b1000111: c <= 9'b100100010;
				8'b1011111: c <= 9'b110001100;
				8'b1110100: c <= 9'b11010100;
				8'b101101: c <= 9'b110000001;
				8'b1010011: c <= 9'b111011100;
				8'b1100001: c <= 9'b110011111;
				8'b110101: c <= 9'b101011;
				8'b1000100: c <= 9'b100001101;
				8'b1010001: c <= 9'b1100100;
				8'b1010100: c <= 9'b1110100;
				8'b1100110: c <= 9'b111111101;
				8'b101010: c <= 9'b110000001;
				8'b1011110: c <= 9'b11101101;
				8'b1100111: c <= 9'b110000;
				8'b1011010: c <= 9'b101101101;
				8'b1000010: c <= 9'b100011111;
				8'b111101: c <= 9'b1000000;
				8'b110000: c <= 9'b1011011;
				8'b111110: c <= 9'b11110011;
				8'b1100010: c <= 9'b11101000;
				8'b1110000: c <= 9'b101100100;
				8'b1101001: c <= 9'b100;
				8'b1110011: c <= 9'b100000101;
				8'b1001100: c <= 9'b101001100;
				8'b100001: c <= 9'b101111001;
				8'b1000110: c <= 9'b1011000;
				8'b1110010: c <= 9'b110000011;
				8'b1010000: c <= 9'b10011011;
				8'b1111010: c <= 9'b10101001;
				8'b1010101: c <= 9'b1101000;
				8'b111011: c <= 9'b11011101;
				8'b1001101: c <= 9'b110010101;
				8'b111111: c <= 9'b11000111;
				8'b1101110: c <= 9'b11001111;
				8'b1111011: c <= 9'b11011110;
				8'b1001011: c <= 9'b11110100;
				8'b1101111: c <= 9'b111011100;
				8'b1101000: c <= 9'b10000000;
				8'b101100: c <= 9'b1001101;
				8'b100100: c <= 9'b1101001;
				8'b1111000: c <= 9'b1010001;
				8'b1000101: c <= 9'b10100;
				8'b1011001: c <= 9'b1111011;
				8'b110100: c <= 9'b111111011;
				8'b1111001: c <= 9'b10000101;
				8'b1110001: c <= 9'b1001101;
				8'b1001111: c <= 9'b11110000;
				8'b1100101: c <= 9'b101001000;
				8'b1111110: c <= 9'b11101001;
				8'b1111100: c <= 9'b10000;
				8'b1010110: c <= 9'b1101010;
				8'b110010: c <= 9'b1010011;
				8'b1101101: c <= 9'b11001110;
				8'b100011: c <= 9'b100;
				8'b1110101: c <= 9'b111110101;
				8'b1111101: c <= 9'b11000100;
				8'b101001: c <= 9'b100010011;
				8'b1010010: c <= 9'b111101001;
				8'b1011000: c <= 9'b11010;
				8'b101110: c <= 9'b10011100;
				8'b1000001: c <= 9'b11100010;
				default: c <= 9'b0;
			endcase
			9'b101100100 : case(di)
				8'b1000011: c <= 9'b1111011;
				8'b101000: c <= 9'b1111110;
				8'b111010: c <= 9'b101011;
				8'b110110: c <= 9'b1100000;
				8'b1100100: c <= 9'b1100011;
				8'b1000000: c <= 9'b10000110;
				8'b1110110: c <= 9'b110100000;
				8'b100101: c <= 9'b100000111;
				8'b101111: c <= 9'b111001110;
				8'b100110: c <= 9'b10010110;
				8'b1100011: c <= 9'b100010101;
				8'b1001000: c <= 9'b10011010;
				8'b111000: c <= 9'b111100000;
				8'b110001: c <= 9'b111001001;
				8'b1010111: c <= 9'b101010010;
				8'b1001110: c <= 9'b101110000;
				8'b1101010: c <= 9'b11101011;
				8'b1001001: c <= 9'b1111111;
				8'b1100000: c <= 9'b110101001;
				8'b110111: c <= 9'b10011001;
				8'b1011101: c <= 9'b1010011;
				8'b1011011: c <= 9'b110011110;
				8'b111001: c <= 9'b111011011;
				8'b1001010: c <= 9'b111001101;
				8'b110011: c <= 9'b101001000;
				8'b1101100: c <= 9'b111101101;
				8'b1110111: c <= 9'b11110100;
				8'b101011: c <= 9'b100101100;
				8'b1101011: c <= 9'b11100011;
				8'b111100: c <= 9'b101011001;
				8'b1000111: c <= 9'b110101010;
				8'b1011111: c <= 9'b1100101;
				8'b1110100: c <= 9'b110100010;
				8'b101101: c <= 9'b101011000;
				8'b1010011: c <= 9'b101110001;
				8'b1100001: c <= 9'b100100010;
				8'b110101: c <= 9'b11110;
				8'b1000100: c <= 9'b111100110;
				8'b1010001: c <= 9'b100101100;
				8'b1010100: c <= 9'b111010001;
				8'b1100110: c <= 9'b110110011;
				8'b101010: c <= 9'b110001100;
				8'b1011110: c <= 9'b101001;
				8'b1100111: c <= 9'b101010010;
				8'b1011010: c <= 9'b11110010;
				8'b1000010: c <= 9'b1111010;
				8'b111101: c <= 9'b10111;
				8'b110000: c <= 9'b110100100;
				8'b111110: c <= 9'b110;
				8'b1100010: c <= 9'b110101011;
				8'b1110000: c <= 9'b100011111;
				8'b1101001: c <= 9'b10001101;
				8'b1110011: c <= 9'b10;
				8'b1001100: c <= 9'b101110101;
				8'b100001: c <= 9'b100000001;
				8'b1000110: c <= 9'b10011000;
				8'b1110010: c <= 9'b111111010;
				8'b1010000: c <= 9'b101101111;
				8'b1111010: c <= 9'b111100;
				8'b1010101: c <= 9'b10000001;
				8'b111011: c <= 9'b100011101;
				8'b1001101: c <= 9'b11100010;
				8'b111111: c <= 9'b111010001;
				8'b1101110: c <= 9'b1001010;
				8'b1111011: c <= 9'b110001111;
				8'b1001011: c <= 9'b10000111;
				8'b1101111: c <= 9'b110111100;
				8'b1101000: c <= 9'b111010110;
				8'b101100: c <= 9'b1000101;
				8'b100100: c <= 9'b11101000;
				8'b1111000: c <= 9'b101011011;
				8'b1000101: c <= 9'b11111011;
				8'b1011001: c <= 9'b100101100;
				8'b110100: c <= 9'b100111110;
				8'b1111001: c <= 9'b110100000;
				8'b1110001: c <= 9'b11110011;
				8'b1001111: c <= 9'b10101000;
				8'b1100101: c <= 9'b101;
				8'b1111110: c <= 9'b1010111;
				8'b1111100: c <= 9'b100011010;
				8'b1010110: c <= 9'b10110;
				8'b110010: c <= 9'b100001001;
				8'b1101101: c <= 9'b10010111;
				8'b100011: c <= 9'b10111001;
				8'b1110101: c <= 9'b1010010;
				8'b1111101: c <= 9'b11010;
				8'b101001: c <= 9'b10101001;
				8'b1010010: c <= 9'b110000111;
				8'b1011000: c <= 9'b110100001;
				8'b101110: c <= 9'b11110011;
				8'b1000001: c <= 9'b1000010;
				default: c <= 9'b0;
			endcase
			9'b10010100 : case(di)
				8'b1000011: c <= 9'b100101001;
				8'b101000: c <= 9'b110101110;
				8'b111010: c <= 9'b11100;
				8'b110110: c <= 9'b10010100;
				8'b1100100: c <= 9'b100000010;
				8'b1000000: c <= 9'b101100;
				8'b1110110: c <= 9'b10001001;
				8'b100101: c <= 9'b1011011;
				8'b101111: c <= 9'b1101101;
				8'b100110: c <= 9'b110001100;
				8'b1100011: c <= 9'b1101010;
				8'b1001000: c <= 9'b110000001;
				8'b111000: c <= 9'b101100011;
				8'b110001: c <= 9'b100010100;
				8'b1010111: c <= 9'b110100000;
				8'b1001110: c <= 9'b1101010;
				8'b1101010: c <= 9'b111100000;
				8'b1001001: c <= 9'b111101101;
				8'b1100000: c <= 9'b10000010;
				8'b110111: c <= 9'b110011;
				8'b1011101: c <= 9'b11111000;
				8'b1011011: c <= 9'b1001100;
				8'b111001: c <= 9'b1000100;
				8'b1001010: c <= 9'b100100010;
				8'b110011: c <= 9'b10011010;
				8'b1101100: c <= 9'b10111110;
				8'b1110111: c <= 9'b110000;
				8'b101011: c <= 9'b100111111;
				8'b1101011: c <= 9'b110010011;
				8'b111100: c <= 9'b11000110;
				8'b1000111: c <= 9'b10111011;
				8'b1011111: c <= 9'b1111010;
				8'b1110100: c <= 9'b101011110;
				8'b101101: c <= 9'b101000110;
				8'b1010011: c <= 9'b101110010;
				8'b1100001: c <= 9'b100010011;
				8'b110101: c <= 9'b110011100;
				8'b1000100: c <= 9'b1100110;
				8'b1010001: c <= 9'b1000;
				8'b1010100: c <= 9'b100010100;
				8'b1100110: c <= 9'b111001001;
				8'b101010: c <= 9'b10110001;
				8'b1011110: c <= 9'b111000;
				8'b1100111: c <= 9'b1110101;
				8'b1011010: c <= 9'b111100010;
				8'b1000010: c <= 9'b101000001;
				8'b111101: c <= 9'b110111011;
				8'b110000: c <= 9'b111101010;
				8'b111110: c <= 9'b1010111;
				8'b1100010: c <= 9'b10000111;
				8'b1110000: c <= 9'b10110101;
				8'b1101001: c <= 9'b111111110;
				8'b1110011: c <= 9'b110111001;
				8'b1001100: c <= 9'b1011;
				8'b100001: c <= 9'b100000001;
				8'b1000110: c <= 9'b1101111;
				8'b1110010: c <= 9'b111100100;
				8'b1010000: c <= 9'b110100;
				8'b1111010: c <= 9'b10111;
				8'b1010101: c <= 9'b1110010;
				8'b111011: c <= 9'b100111110;
				8'b1001101: c <= 9'b101111110;
				8'b111111: c <= 9'b111001010;
				8'b1101110: c <= 9'b101010;
				8'b1111011: c <= 9'b10110010;
				8'b1001011: c <= 9'b100010000;
				8'b1101111: c <= 9'b1010000;
				8'b1101000: c <= 9'b111001011;
				8'b101100: c <= 9'b10001010;
				8'b100100: c <= 9'b1010110;
				8'b1111000: c <= 9'b111101010;
				8'b1000101: c <= 9'b10110011;
				8'b1011001: c <= 9'b11001011;
				8'b110100: c <= 9'b101100000;
				8'b1111001: c <= 9'b100010;
				8'b1110001: c <= 9'b100101;
				8'b1001111: c <= 9'b111000;
				8'b1100101: c <= 9'b1;
				8'b1111110: c <= 9'b100100110;
				8'b1111100: c <= 9'b11111101;
				8'b1010110: c <= 9'b10111110;
				8'b110010: c <= 9'b111111000;
				8'b1101101: c <= 9'b110001010;
				8'b100011: c <= 9'b1111100;
				8'b1110101: c <= 9'b11100101;
				8'b1111101: c <= 9'b1010001;
				8'b101001: c <= 9'b101001100;
				8'b1010010: c <= 9'b100101001;
				8'b1011000: c <= 9'b1100010;
				8'b101110: c <= 9'b10001010;
				8'b1000001: c <= 9'b111010001;
				default: c <= 9'b0;
			endcase
			9'b101110 : case(di)
				8'b1000011: c <= 9'b10010001;
				8'b101000: c <= 9'b111010111;
				8'b111010: c <= 9'b1111111;
				8'b110110: c <= 9'b1111101;
				8'b1100100: c <= 9'b1111010;
				8'b1000000: c <= 9'b100011;
				8'b1110110: c <= 9'b100001110;
				8'b100101: c <= 9'b101001;
				8'b101111: c <= 9'b110011100;
				8'b100110: c <= 9'b100100;
				8'b1100011: c <= 9'b110010100;
				8'b1001000: c <= 9'b101111010;
				8'b111000: c <= 9'b101111001;
				8'b110001: c <= 9'b11101001;
				8'b1010111: c <= 9'b111010010;
				8'b1001110: c <= 9'b1001101;
				8'b1101010: c <= 9'b101100110;
				8'b1001001: c <= 9'b110110000;
				8'b1100000: c <= 9'b101000;
				8'b110111: c <= 9'b1000000;
				8'b1011101: c <= 9'b10111101;
				8'b1011011: c <= 9'b101000101;
				8'b111001: c <= 9'b111101;
				8'b1001010: c <= 9'b10110110;
				8'b110011: c <= 9'b1110;
				8'b1101100: c <= 9'b10001100;
				8'b1110111: c <= 9'b111011111;
				8'b101011: c <= 9'b110001100;
				8'b1101011: c <= 9'b11001011;
				8'b111100: c <= 9'b1101111;
				8'b1000111: c <= 9'b1111;
				8'b1011111: c <= 9'b111010001;
				8'b1110100: c <= 9'b11011011;
				8'b101101: c <= 9'b1100001;
				8'b1010011: c <= 9'b1000100;
				8'b1100001: c <= 9'b111001100;
				8'b110101: c <= 9'b11100010;
				8'b1000100: c <= 9'b11011001;
				8'b1010001: c <= 9'b1110001;
				8'b1010100: c <= 9'b101101010;
				8'b1100110: c <= 9'b10111111;
				8'b101010: c <= 9'b100001010;
				8'b1011110: c <= 9'b100101110;
				8'b1100111: c <= 9'b11010101;
				8'b1011010: c <= 9'b1110001;
				8'b1000010: c <= 9'b111000111;
				8'b111101: c <= 9'b1111001;
				8'b110000: c <= 9'b101000010;
				8'b111110: c <= 9'b1000;
				8'b1100010: c <= 9'b10011000;
				8'b1110000: c <= 9'b111101100;
				8'b1101001: c <= 9'b1011110;
				8'b1110011: c <= 9'b1101111;
				8'b1001100: c <= 9'b111011011;
				8'b100001: c <= 9'b101001000;
				8'b1000110: c <= 9'b100110;
				8'b1110010: c <= 9'b1011111;
				8'b1010000: c <= 9'b1001011;
				8'b1111010: c <= 9'b110100100;
				8'b1010101: c <= 9'b11110111;
				8'b111011: c <= 9'b100001001;
				8'b1001101: c <= 9'b101011101;
				8'b111111: c <= 9'b111101111;
				8'b1101110: c <= 9'b110111110;
				8'b1111011: c <= 9'b100101110;
				8'b1001011: c <= 9'b101100101;
				8'b1101111: c <= 9'b100010101;
				8'b1101000: c <= 9'b111111101;
				8'b101100: c <= 9'b1000111;
				8'b100100: c <= 9'b101111000;
				8'b1111000: c <= 9'b1001;
				8'b1000101: c <= 9'b100111011;
				8'b1011001: c <= 9'b11110000;
				8'b110100: c <= 9'b1011110;
				8'b1111001: c <= 9'b110001110;
				8'b1110001: c <= 9'b1101010;
				8'b1001111: c <= 9'b11100001;
				8'b1100101: c <= 9'b111110101;
				8'b1111110: c <= 9'b101100100;
				8'b1111100: c <= 9'b10101011;
				8'b1010110: c <= 9'b11100;
				8'b110010: c <= 9'b10000010;
				8'b1101101: c <= 9'b10110111;
				8'b100011: c <= 9'b10000;
				8'b1110101: c <= 9'b1011001;
				8'b1111101: c <= 9'b11001010;
				8'b101001: c <= 9'b10011001;
				8'b1010010: c <= 9'b1000;
				8'b1011000: c <= 9'b111100000;
				8'b101110: c <= 9'b101001001;
				8'b1000001: c <= 9'b111111010;
				default: c <= 9'b0;
			endcase
			9'b1110 : case(di)
				8'b1000011: c <= 9'b10000011;
				8'b101000: c <= 9'b110110000;
				8'b111010: c <= 9'b111000;
				8'b110110: c <= 9'b10000001;
				8'b1100100: c <= 9'b100100011;
				8'b1000000: c <= 9'b11001;
				8'b1110110: c <= 9'b110111;
				8'b100101: c <= 9'b111110101;
				8'b101111: c <= 9'b100010110;
				8'b100110: c <= 9'b10011101;
				8'b1100011: c <= 9'b11110110;
				8'b1001000: c <= 9'b111000011;
				8'b111000: c <= 9'b100100;
				8'b110001: c <= 9'b1110011;
				8'b1010111: c <= 9'b111100;
				8'b1001110: c <= 9'b110001000;
				8'b1101010: c <= 9'b11;
				8'b1001001: c <= 9'b11110111;
				8'b1100000: c <= 9'b11001001;
				8'b110111: c <= 9'b1101000;
				8'b1011101: c <= 9'b10110010;
				8'b1011011: c <= 9'b100111100;
				8'b111001: c <= 9'b101100110;
				8'b1001010: c <= 9'b111010110;
				8'b110011: c <= 9'b1001000;
				8'b1101100: c <= 9'b110;
				8'b1110111: c <= 9'b11000010;
				8'b101011: c <= 9'b111111001;
				8'b1101011: c <= 9'b100111100;
				8'b111100: c <= 9'b11011010;
				8'b1000111: c <= 9'b11011001;
				8'b1011111: c <= 9'b110110100;
				8'b1110100: c <= 9'b1100010;
				8'b101101: c <= 9'b111011011;
				8'b1010011: c <= 9'b11011011;
				8'b1100001: c <= 9'b1011111;
				8'b110101: c <= 9'b11110111;
				8'b1000100: c <= 9'b110101011;
				8'b1010001: c <= 9'b100000100;
				8'b1010100: c <= 9'b111100000;
				8'b1100110: c <= 9'b100101111;
				8'b101010: c <= 9'b1100110;
				8'b1011110: c <= 9'b10000011;
				8'b1100111: c <= 9'b110000;
				8'b1011010: c <= 9'b11110;
				8'b1000010: c <= 9'b100010010;
				8'b111101: c <= 9'b100101010;
				8'b110000: c <= 9'b100001111;
				8'b111110: c <= 9'b11001001;
				8'b1100010: c <= 9'b101010101;
				8'b1110000: c <= 9'b100011100;
				8'b1101001: c <= 9'b100001;
				8'b1110011: c <= 9'b111100101;
				8'b1001100: c <= 9'b101101000;
				8'b100001: c <= 9'b11011101;
				8'b1000110: c <= 9'b10111101;
				8'b1110010: c <= 9'b101010110;
				8'b1010000: c <= 9'b111101;
				8'b1111010: c <= 9'b110000011;
				8'b1010101: c <= 9'b111100001;
				8'b111011: c <= 9'b111100000;
				8'b1001101: c <= 9'b1111010;
				8'b111111: c <= 9'b111011101;
				8'b1101110: c <= 9'b100010101;
				8'b1111011: c <= 9'b100001111;
				8'b1001011: c <= 9'b111101010;
				8'b1101111: c <= 9'b111100111;
				8'b1101000: c <= 9'b111000;
				8'b101100: c <= 9'b110111110;
				8'b100100: c <= 9'b111110001;
				8'b1111000: c <= 9'b100000101;
				8'b1000101: c <= 9'b100010;
				8'b1011001: c <= 9'b111100000;
				8'b110100: c <= 9'b101011110;
				8'b1111001: c <= 9'b11000100;
				8'b1110001: c <= 9'b101100110;
				8'b1001111: c <= 9'b10101100;
				8'b1100101: c <= 9'b1001011;
				8'b1111110: c <= 9'b100111111;
				8'b1111100: c <= 9'b11010010;
				8'b1010110: c <= 9'b1;
				8'b110010: c <= 9'b1111000;
				8'b1101101: c <= 9'b10111110;
				8'b100011: c <= 9'b1000110;
				8'b1110101: c <= 9'b111011010;
				8'b1111101: c <= 9'b10001100;
				8'b101001: c <= 9'b101111010;
				8'b1010010: c <= 9'b110110010;
				8'b1011000: c <= 9'b110100010;
				8'b101110: c <= 9'b10111100;
				8'b1000001: c <= 9'b110100111;
				default: c <= 9'b0;
			endcase
			9'b1 : case(di)
				8'b1000011: c <= 9'b100111010;
				8'b101000: c <= 9'b11110100;
				8'b111010: c <= 9'b10100011;
				8'b110110: c <= 9'b111001100;
				8'b1100100: c <= 9'b101010101;
				8'b1000000: c <= 9'b1001101;
				8'b1110110: c <= 9'b101100110;
				8'b100101: c <= 9'b10110001;
				8'b101111: c <= 9'b100111111;
				8'b100110: c <= 9'b1001100;
				8'b1100011: c <= 9'b100000111;
				8'b1001000: c <= 9'b1110100;
				8'b111000: c <= 9'b111101;
				8'b110001: c <= 9'b100001101;
				8'b1010111: c <= 9'b110110110;
				8'b1001110: c <= 9'b101000101;
				8'b1101010: c <= 9'b101001001;
				8'b1001001: c <= 9'b11010111;
				8'b1100000: c <= 9'b10000110;
				8'b110111: c <= 9'b100011011;
				8'b1011101: c <= 9'b10001101;
				8'b1011011: c <= 9'b11001001;
				8'b111001: c <= 9'b1001111;
				8'b1001010: c <= 9'b10111001;
				8'b110011: c <= 9'b101110000;
				8'b1101100: c <= 9'b11011101;
				8'b1110111: c <= 9'b1011111;
				8'b101011: c <= 9'b110000101;
				8'b1101011: c <= 9'b11110100;
				8'b111100: c <= 9'b110000000;
				8'b1000111: c <= 9'b100111001;
				8'b1011111: c <= 9'b1100011;
				8'b1110100: c <= 9'b101011101;
				8'b101101: c <= 9'b11011001;
				8'b1010011: c <= 9'b1000;
				8'b1100001: c <= 9'b10000101;
				8'b110101: c <= 9'b10011010;
				8'b1000100: c <= 9'b1001101;
				8'b1010001: c <= 9'b100100110;
				8'b1010100: c <= 9'b11110110;
				8'b1100110: c <= 9'b11110011;
				8'b101010: c <= 9'b101100101;
				8'b1011110: c <= 9'b101001;
				8'b1100111: c <= 9'b10110111;
				8'b1011010: c <= 9'b1011100;
				8'b1000010: c <= 9'b11110101;
				8'b111101: c <= 9'b1010111;
				8'b110000: c <= 9'b111100011;
				8'b111110: c <= 9'b100010001;
				8'b1100010: c <= 9'b110101;
				8'b1110000: c <= 9'b110001011;
				8'b1101001: c <= 9'b100100110;
				8'b1110011: c <= 9'b100101111;
				8'b1001100: c <= 9'b111100110;
				8'b100001: c <= 9'b10010101;
				8'b1000110: c <= 9'b10011000;
				8'b1110010: c <= 9'b1111101;
				8'b1010000: c <= 9'b111110110;
				8'b1111010: c <= 9'b1011010;
				8'b1010101: c <= 9'b101100111;
				8'b111011: c <= 9'b100010111;
				8'b1001101: c <= 9'b1100011;
				8'b111111: c <= 9'b111000111;
				8'b1101110: c <= 9'b110010010;
				8'b1111011: c <= 9'b111011110;
				8'b1001011: c <= 9'b1011000;
				8'b1101111: c <= 9'b111111111;
				8'b1101000: c <= 9'b110000011;
				8'b101100: c <= 9'b101011010;
				8'b100100: c <= 9'b10101000;
				8'b1111000: c <= 9'b110111001;
				8'b1000101: c <= 9'b101001001;
				8'b1011001: c <= 9'b10110001;
				8'b110100: c <= 9'b1110100;
				8'b1111001: c <= 9'b111100;
				8'b1110001: c <= 9'b110110111;
				8'b1001111: c <= 9'b11010011;
				8'b1100101: c <= 9'b101011110;
				8'b1111110: c <= 9'b110100011;
				8'b1111100: c <= 9'b11110101;
				8'b1010110: c <= 9'b100011101;
				8'b110010: c <= 9'b1001101;
				8'b1101101: c <= 9'b111010000;
				8'b100011: c <= 9'b10101001;
				8'b1110101: c <= 9'b101100011;
				8'b1111101: c <= 9'b11100100;
				8'b101001: c <= 9'b111111111;
				8'b1010010: c <= 9'b101001001;
				8'b1011000: c <= 9'b100000101;
				8'b101110: c <= 9'b10001101;
				8'b1000001: c <= 9'b1111110;
				default: c <= 9'b0;
			endcase
			9'b111000100 : case(di)
				8'b1000011: c <= 9'b110001000;
				8'b101000: c <= 9'b10100011;
				8'b111010: c <= 9'b110001000;
				8'b110110: c <= 9'b11001001;
				8'b1100100: c <= 9'b100000010;
				8'b1000000: c <= 9'b10111011;
				8'b1110110: c <= 9'b100;
				8'b100101: c <= 9'b100000000;
				8'b101111: c <= 9'b110011111;
				8'b100110: c <= 9'b1101010;
				8'b1100011: c <= 9'b101101110;
				8'b1001000: c <= 9'b110111010;
				8'b111000: c <= 9'b10100;
				8'b110001: c <= 9'b111100000;
				8'b1010111: c <= 9'b111110110;
				8'b1001110: c <= 9'b111001010;
				8'b1101010: c <= 9'b10001000;
				8'b1001001: c <= 9'b110001;
				8'b1100000: c <= 9'b10000;
				8'b110111: c <= 9'b10011111;
				8'b1011101: c <= 9'b11001011;
				8'b1011011: c <= 9'b101110010;
				8'b111001: c <= 9'b11010101;
				8'b1001010: c <= 9'b101100001;
				8'b110011: c <= 9'b10111101;
				8'b1101100: c <= 9'b100010110;
				8'b1110111: c <= 9'b101111001;
				8'b101011: c <= 9'b110001110;
				8'b1101011: c <= 9'b101100;
				8'b111100: c <= 9'b111110011;
				8'b1000111: c <= 9'b110011;
				8'b1011111: c <= 9'b111101010;
				8'b1110100: c <= 9'b110011110;
				8'b101101: c <= 9'b1110001;
				8'b1010011: c <= 9'b10111100;
				8'b1100001: c <= 9'b100001111;
				8'b110101: c <= 9'b110100010;
				8'b1000100: c <= 9'b111001110;
				8'b1010001: c <= 9'b111111001;
				8'b1010100: c <= 9'b111101100;
				8'b1100110: c <= 9'b100001;
				8'b101010: c <= 9'b11111000;
				8'b1011110: c <= 9'b111011100;
				8'b1100111: c <= 9'b110111;
				8'b1011010: c <= 9'b10111110;
				8'b1000010: c <= 9'b1101000;
				8'b111101: c <= 9'b110101010;
				8'b110000: c <= 9'b10111000;
				8'b111110: c <= 9'b11100010;
				8'b1100010: c <= 9'b11001011;
				8'b1110000: c <= 9'b110101100;
				8'b1101001: c <= 9'b11111001;
				8'b1110011: c <= 9'b100001001;
				8'b1001100: c <= 9'b100111100;
				8'b100001: c <= 9'b100101001;
				8'b1000110: c <= 9'b1111000;
				8'b1110010: c <= 9'b11011000;
				8'b1010000: c <= 9'b110000011;
				8'b1111010: c <= 9'b101001;
				8'b1010101: c <= 9'b1010001;
				8'b111011: c <= 9'b11110110;
				8'b1001101: c <= 9'b10011;
				8'b111111: c <= 9'b10110;
				8'b1101110: c <= 9'b1101111;
				8'b1111011: c <= 9'b11100;
				8'b1001011: c <= 9'b100100011;
				8'b1101111: c <= 9'b110011111;
				8'b1101000: c <= 9'b10111001;
				8'b101100: c <= 9'b111100000;
				8'b100100: c <= 9'b100100010;
				8'b1111000: c <= 9'b1011011;
				8'b1000101: c <= 9'b111000110;
				8'b1011001: c <= 9'b1011001;
				8'b110100: c <= 9'b100001;
				8'b1111001: c <= 9'b101110100;
				8'b1110001: c <= 9'b110100011;
				8'b1001111: c <= 9'b1;
				8'b1100101: c <= 9'b111111001;
				8'b1111110: c <= 9'b11001011;
				8'b1111100: c <= 9'b1100110;
				8'b1010110: c <= 9'b10010101;
				8'b110010: c <= 9'b1010110;
				8'b1101101: c <= 9'b110100101;
				8'b100011: c <= 9'b10111111;
				8'b1110101: c <= 9'b10101011;
				8'b1111101: c <= 9'b101110111;
				8'b101001: c <= 9'b100110110;
				8'b1010010: c <= 9'b101101101;
				8'b1011000: c <= 9'b100010011;
				8'b101110: c <= 9'b1110010;
				8'b1000001: c <= 9'b11101111;
				default: c <= 9'b0;
			endcase
			9'b111111101 : case(di)
				8'b1000011: c <= 9'b110000001;
				8'b101000: c <= 9'b1001101;
				8'b111010: c <= 9'b100110100;
				8'b110110: c <= 9'b100000010;
				8'b1100100: c <= 9'b11001111;
				8'b1000000: c <= 9'b10101011;
				8'b1110110: c <= 9'b100011000;
				8'b100101: c <= 9'b11110101;
				8'b101111: c <= 9'b111110101;
				8'b100110: c <= 9'b101101001;
				8'b1100011: c <= 9'b111001111;
				8'b1001000: c <= 9'b111011100;
				8'b111000: c <= 9'b110001110;
				8'b110001: c <= 9'b11110000;
				8'b1010111: c <= 9'b10110;
				8'b1001110: c <= 9'b10111110;
				8'b1101010: c <= 9'b101000011;
				8'b1001001: c <= 9'b110111001;
				8'b1100000: c <= 9'b1100100;
				8'b110111: c <= 9'b100011100;
				8'b1011101: c <= 9'b110010;
				8'b1011011: c <= 9'b1110111;
				8'b111001: c <= 9'b111110110;
				8'b1001010: c <= 9'b11010101;
				8'b110011: c <= 9'b101000111;
				8'b1101100: c <= 9'b101110011;
				8'b1110111: c <= 9'b10000010;
				8'b101011: c <= 9'b11101011;
				8'b1101011: c <= 9'b100010100;
				8'b111100: c <= 9'b101111010;
				8'b1000111: c <= 9'b11001;
				8'b1011111: c <= 9'b110111001;
				8'b1110100: c <= 9'b101001000;
				8'b101101: c <= 9'b11111010;
				8'b1010011: c <= 9'b1001001;
				8'b1100001: c <= 9'b1000001;
				8'b110101: c <= 9'b110010010;
				8'b1000100: c <= 9'b101101111;
				8'b1010001: c <= 9'b11011110;
				8'b1010100: c <= 9'b10101010;
				8'b1100110: c <= 9'b101011101;
				8'b101010: c <= 9'b101110100;
				8'b1011110: c <= 9'b111010100;
				8'b1100111: c <= 9'b101100110;
				8'b1011010: c <= 9'b11011011;
				8'b1000010: c <= 9'b110101111;
				8'b111101: c <= 9'b110101;
				8'b110000: c <= 9'b11000111;
				8'b111110: c <= 9'b11010010;
				8'b1100010: c <= 9'b1000001;
				8'b1110000: c <= 9'b110010110;
				8'b1101001: c <= 9'b110110110;
				8'b1110011: c <= 9'b11111110;
				8'b1001100: c <= 9'b10010101;
				8'b100001: c <= 9'b1010111;
				8'b1000110: c <= 9'b11110010;
				8'b1110010: c <= 9'b101;
				8'b1010000: c <= 9'b100010;
				8'b1111010: c <= 9'b1101111;
				8'b1010101: c <= 9'b111110110;
				8'b111011: c <= 9'b100000001;
				8'b1001101: c <= 9'b110100;
				8'b111111: c <= 9'b111100111;
				8'b1101110: c <= 9'b10011;
				8'b1111011: c <= 9'b101100110;
				8'b1001011: c <= 9'b11111101;
				8'b1101111: c <= 9'b111000111;
				8'b1101000: c <= 9'b111000110;
				8'b101100: c <= 9'b111101100;
				8'b100100: c <= 9'b1110011;
				8'b1111000: c <= 9'b10000000;
				8'b1000101: c <= 9'b10111100;
				8'b1011001: c <= 9'b11011011;
				8'b110100: c <= 9'b11100100;
				8'b1111001: c <= 9'b110010010;
				8'b1110001: c <= 9'b111101001;
				8'b1001111: c <= 9'b101100111;
				8'b1100101: c <= 9'b111110110;
				8'b1111110: c <= 9'b100001111;
				8'b1111100: c <= 9'b1001111;
				8'b1010110: c <= 9'b100101111;
				8'b110010: c <= 9'b110101010;
				8'b1101101: c <= 9'b1000010;
				8'b100011: c <= 9'b11110100;
				8'b1110101: c <= 9'b11001011;
				8'b1111101: c <= 9'b101100000;
				8'b101001: c <= 9'b10111010;
				8'b1010010: c <= 9'b11000000;
				8'b1011000: c <= 9'b110100111;
				8'b101110: c <= 9'b100111111;
				8'b1000001: c <= 9'b110101110;
				default: c <= 9'b0;
			endcase
			9'b1000010 : case(di)
				8'b1000011: c <= 9'b110011;
				8'b101000: c <= 9'b110101100;
				8'b111010: c <= 9'b100000000;
				8'b110110: c <= 9'b111101;
				8'b1100100: c <= 9'b100001101;
				8'b1000000: c <= 9'b111100111;
				8'b1110110: c <= 9'b110000010;
				8'b100101: c <= 9'b111011010;
				8'b101111: c <= 9'b110001111;
				8'b100110: c <= 9'b101101001;
				8'b1100011: c <= 9'b101110011;
				8'b1001000: c <= 9'b110110010;
				8'b111000: c <= 9'b110100010;
				8'b110001: c <= 9'b11000;
				8'b1010111: c <= 9'b1000010;
				8'b1001110: c <= 9'b110001001;
				8'b1101010: c <= 9'b101011101;
				8'b1001001: c <= 9'b100011;
				8'b1100000: c <= 9'b11111101;
				8'b110111: c <= 9'b110110110;
				8'b1011101: c <= 9'b110000011;
				8'b1011011: c <= 9'b110010110;
				8'b111001: c <= 9'b1100101;
				8'b1001010: c <= 9'b111100111;
				8'b110011: c <= 9'b100101101;
				8'b1101100: c <= 9'b1111010;
				8'b1110111: c <= 9'b11000110;
				8'b101011: c <= 9'b1100000;
				8'b1101011: c <= 9'b100111111;
				8'b111100: c <= 9'b11001110;
				8'b1000111: c <= 9'b1100000;
				8'b1011111: c <= 9'b101100010;
				8'b1110100: c <= 9'b100111100;
				8'b101101: c <= 9'b1110000;
				8'b1010011: c <= 9'b1100;
				8'b1100001: c <= 9'b100110100;
				8'b110101: c <= 9'b11100101;
				8'b1000100: c <= 9'b11111100;
				8'b1010001: c <= 9'b1110010;
				8'b1010100: c <= 9'b110100101;
				8'b1100110: c <= 9'b101100011;
				8'b101010: c <= 9'b111101111;
				8'b1011110: c <= 9'b110011010;
				8'b1100111: c <= 9'b10010011;
				8'b1011010: c <= 9'b110100010;
				8'b1000010: c <= 9'b1101110;
				8'b111101: c <= 9'b101101001;
				8'b110000: c <= 9'b111010000;
				8'b111110: c <= 9'b111010001;
				8'b1100010: c <= 9'b10010001;
				8'b1110000: c <= 9'b10000111;
				8'b1101001: c <= 9'b11110;
				8'b1110011: c <= 9'b11000110;
				8'b1001100: c <= 9'b110101;
				8'b100001: c <= 9'b101000010;
				8'b1000110: c <= 9'b10010;
				8'b1110010: c <= 9'b11101011;
				8'b1010000: c <= 9'b101100110;
				8'b1111010: c <= 9'b110001011;
				8'b1010101: c <= 9'b10000010;
				8'b111011: c <= 9'b111101111;
				8'b1001101: c <= 9'b1110010;
				8'b111111: c <= 9'b110100;
				8'b1101110: c <= 9'b11000001;
				8'b1111011: c <= 9'b111111101;
				8'b1001011: c <= 9'b100111011;
				8'b1101111: c <= 9'b10111100;
				8'b1101000: c <= 9'b10100111;
				8'b101100: c <= 9'b101100110;
				8'b100100: c <= 9'b111111101;
				8'b1111000: c <= 9'b10000111;
				8'b1000101: c <= 9'b111011110;
				8'b1011001: c <= 9'b11111001;
				8'b110100: c <= 9'b1110111;
				8'b1111001: c <= 9'b101000110;
				8'b1110001: c <= 9'b11100100;
				8'b1001111: c <= 9'b1110010;
				8'b1100101: c <= 9'b11001000;
				8'b1111110: c <= 9'b1101;
				8'b1111100: c <= 9'b111101110;
				8'b1010110: c <= 9'b11111001;
				8'b110010: c <= 9'b1000;
				8'b1101101: c <= 9'b1100110;
				8'b100011: c <= 9'b111100011;
				8'b1110101: c <= 9'b110011000;
				8'b1111101: c <= 9'b111110101;
				8'b101001: c <= 9'b110110010;
				8'b1010010: c <= 9'b111111010;
				8'b1011000: c <= 9'b1011010;
				8'b101110: c <= 9'b101111010;
				8'b1000001: c <= 9'b1110001;
				default: c <= 9'b0;
			endcase
			9'b101001010 : case(di)
				8'b1000011: c <= 9'b10010;
				8'b101000: c <= 9'b1000;
				8'b111010: c <= 9'b110110010;
				8'b110110: c <= 9'b100011000;
				8'b1100100: c <= 9'b110110;
				8'b1000000: c <= 9'b110011100;
				8'b1110110: c <= 9'b101010001;
				8'b100101: c <= 9'b10100100;
				8'b101111: c <= 9'b100110111;
				8'b100110: c <= 9'b11100101;
				8'b1100011: c <= 9'b10000001;
				8'b1001000: c <= 9'b11000000;
				8'b111000: c <= 9'b11100;
				8'b110001: c <= 9'b10100;
				8'b1010111: c <= 9'b100000001;
				8'b1001110: c <= 9'b10001011;
				8'b1101010: c <= 9'b11001010;
				8'b1001001: c <= 9'b111000;
				8'b1100000: c <= 9'b100111;
				8'b110111: c <= 9'b1000;
				8'b1011101: c <= 9'b101001110;
				8'b1011011: c <= 9'b111101110;
				8'b111001: c <= 9'b1001110;
				8'b1001010: c <= 9'b100010011;
				8'b110011: c <= 9'b11000001;
				8'b1101100: c <= 9'b100110010;
				8'b1110111: c <= 9'b11010001;
				8'b101011: c <= 9'b10011011;
				8'b1101011: c <= 9'b111110101;
				8'b111100: c <= 9'b111000111;
				8'b1000111: c <= 9'b101000110;
				8'b1011111: c <= 9'b10110011;
				8'b1110100: c <= 9'b110010101;
				8'b101101: c <= 9'b111101;
				8'b1010011: c <= 9'b11010100;
				8'b1100001: c <= 9'b101000001;
				8'b110101: c <= 9'b1011;
				8'b1000100: c <= 9'b110110111;
				8'b1010001: c <= 9'b10;
				8'b1010100: c <= 9'b111111010;
				8'b1100110: c <= 9'b110110110;
				8'b101010: c <= 9'b101100110;
				8'b1011110: c <= 9'b110110000;
				8'b1100111: c <= 9'b100010101;
				8'b1011010: c <= 9'b1111110;
				8'b1000010: c <= 9'b110100010;
				8'b111101: c <= 9'b110;
				8'b110000: c <= 9'b100101111;
				8'b111110: c <= 9'b101101;
				8'b1100010: c <= 9'b101101111;
				8'b1110000: c <= 9'b100001010;
				8'b1101001: c <= 9'b100000101;
				8'b1110011: c <= 9'b1000000;
				8'b1001100: c <= 9'b101000011;
				8'b100001: c <= 9'b101101000;
				8'b1000110: c <= 9'b110111000;
				8'b1110010: c <= 9'b100000101;
				8'b1010000: c <= 9'b101000001;
				8'b1111010: c <= 9'b101001111;
				8'b1010101: c <= 9'b110101101;
				8'b111011: c <= 9'b1111111;
				8'b1001101: c <= 9'b110011101;
				8'b111111: c <= 9'b10111101;
				8'b1101110: c <= 9'b1000001;
				8'b1111011: c <= 9'b10110101;
				8'b1001011: c <= 9'b1000010;
				8'b1101111: c <= 9'b10100101;
				8'b1101000: c <= 9'b101010100;
				8'b101100: c <= 9'b100011101;
				8'b100100: c <= 9'b11100010;
				8'b1111000: c <= 9'b101111001;
				8'b1000101: c <= 9'b101001001;
				8'b1011001: c <= 9'b101101;
				8'b110100: c <= 9'b110110100;
				8'b1111001: c <= 9'b101111000;
				8'b1110001: c <= 9'b110001010;
				8'b1001111: c <= 9'b10010;
				8'b1100101: c <= 9'b10011;
				8'b1111110: c <= 9'b11111001;
				8'b1111100: c <= 9'b10001110;
				8'b1010110: c <= 9'b11010001;
				8'b110010: c <= 9'b111001;
				8'b1101101: c <= 9'b10001111;
				8'b100011: c <= 9'b100101011;
				8'b1110101: c <= 9'b11000010;
				8'b1111101: c <= 9'b10111100;
				8'b101001: c <= 9'b11001110;
				8'b1010010: c <= 9'b101001111;
				8'b1011000: c <= 9'b1110111;
				8'b101110: c <= 9'b110101;
				8'b1000001: c <= 9'b100011111;
				default: c <= 9'b0;
			endcase
			9'b1000100 : case(di)
				8'b1000011: c <= 9'b110100000;
				8'b101000: c <= 9'b10111111;
				8'b111010: c <= 9'b101101010;
				8'b110110: c <= 9'b110011101;
				8'b1100100: c <= 9'b111100011;
				8'b1000000: c <= 9'b10111011;
				8'b1110110: c <= 9'b10101111;
				8'b100101: c <= 9'b111101110;
				8'b101111: c <= 9'b111010110;
				8'b100110: c <= 9'b110100111;
				8'b1100011: c <= 9'b111110110;
				8'b1001000: c <= 9'b11100111;
				8'b111000: c <= 9'b111010;
				8'b110001: c <= 9'b110010;
				8'b1010111: c <= 9'b110110100;
				8'b1001110: c <= 9'b110011011;
				8'b1101010: c <= 9'b110011;
				8'b1001001: c <= 9'b101010101;
				8'b1100000: c <= 9'b110000101;
				8'b110111: c <= 9'b110110101;
				8'b1011101: c <= 9'b111000100;
				8'b1011011: c <= 9'b111110011;
				8'b111001: c <= 9'b100011001;
				8'b1001010: c <= 9'b110011101;
				8'b110011: c <= 9'b100101010;
				8'b1101100: c <= 9'b110100000;
				8'b1110111: c <= 9'b10101001;
				8'b101011: c <= 9'b110010111;
				8'b1101011: c <= 9'b100001110;
				8'b111100: c <= 9'b1110010;
				8'b1000111: c <= 9'b1100111;
				8'b1011111: c <= 9'b1001101;
				8'b1110100: c <= 9'b101101;
				8'b101101: c <= 9'b100000010;
				8'b1010011: c <= 9'b110111011;
				8'b1100001: c <= 9'b101101111;
				8'b110101: c <= 9'b100011010;
				8'b1000100: c <= 9'b10000001;
				8'b1010001: c <= 9'b10101000;
				8'b1010100: c <= 9'b1011011;
				8'b1100110: c <= 9'b110111110;
				8'b101010: c <= 9'b101101110;
				8'b1011110: c <= 9'b101111001;
				8'b1100111: c <= 9'b100110011;
				8'b1011010: c <= 9'b1100110;
				8'b1000010: c <= 9'b100000101;
				8'b111101: c <= 9'b110101110;
				8'b110000: c <= 9'b100001110;
				8'b111110: c <= 9'b110111111;
				8'b1100010: c <= 9'b10001000;
				8'b1110000: c <= 9'b1101010;
				8'b1101001: c <= 9'b101000;
				8'b1110011: c <= 9'b11011100;
				8'b1001100: c <= 9'b100101011;
				8'b100001: c <= 9'b110100000;
				8'b1000110: c <= 9'b10100110;
				8'b1110010: c <= 9'b1101100;
				8'b1010000: c <= 9'b1011100;
				8'b1111010: c <= 9'b110010001;
				8'b1010101: c <= 9'b10100110;
				8'b111011: c <= 9'b100011101;
				8'b1001101: c <= 9'b11000111;
				8'b111111: c <= 9'b110100000;
				8'b1101110: c <= 9'b10101100;
				8'b1111011: c <= 9'b111001000;
				8'b1001011: c <= 9'b101010101;
				8'b1101111: c <= 9'b111010000;
				8'b1101000: c <= 9'b10010;
				8'b101100: c <= 9'b111100010;
				8'b100100: c <= 9'b110100000;
				8'b1111000: c <= 9'b100000100;
				8'b1000101: c <= 9'b11011101;
				8'b1011001: c <= 9'b101000;
				8'b110100: c <= 9'b111110000;
				8'b1111001: c <= 9'b110010100;
				8'b1110001: c <= 9'b11110010;
				8'b1001111: c <= 9'b10001001;
				8'b1100101: c <= 9'b111000000;
				8'b1111110: c <= 9'b1100010;
				8'b1111100: c <= 9'b110100000;
				8'b1010110: c <= 9'b110111111;
				8'b110010: c <= 9'b110011100;
				8'b1101101: c <= 9'b10111111;
				8'b100011: c <= 9'b10100011;
				8'b1110101: c <= 9'b11100;
				8'b1111101: c <= 9'b1011010;
				8'b101001: c <= 9'b110011101;
				8'b1010010: c <= 9'b100001011;
				8'b1011000: c <= 9'b110100;
				8'b101110: c <= 9'b11001111;
				8'b1000001: c <= 9'b100100001;
				default: c <= 9'b0;
			endcase
			9'b11110 : case(di)
				8'b1000011: c <= 9'b100000110;
				8'b101000: c <= 9'b111101111;
				8'b111010: c <= 9'b11100000;
				8'b110110: c <= 9'b101011000;
				8'b1100100: c <= 9'b100111100;
				8'b1000000: c <= 9'b110111001;
				8'b1110110: c <= 9'b111011111;
				8'b100101: c <= 9'b101110011;
				8'b101111: c <= 9'b100000010;
				8'b100110: c <= 9'b1010010;
				8'b1100011: c <= 9'b111000101;
				8'b1001000: c <= 9'b111011101;
				8'b111000: c <= 9'b111001111;
				8'b110001: c <= 9'b101011;
				8'b1010111: c <= 9'b110010010;
				8'b1001110: c <= 9'b100001001;
				8'b1101010: c <= 9'b111001000;
				8'b1001001: c <= 9'b11000110;
				8'b1100000: c <= 9'b110101;
				8'b110111: c <= 9'b1111100;
				8'b1011101: c <= 9'b100100111;
				8'b1011011: c <= 9'b111011010;
				8'b111001: c <= 9'b10101;
				8'b1001010: c <= 9'b1100100;
				8'b110011: c <= 9'b11101101;
				8'b1101100: c <= 9'b10001001;
				8'b1110111: c <= 9'b110001101;
				8'b101011: c <= 9'b110101;
				8'b1101011: c <= 9'b11000000;
				8'b111100: c <= 9'b1001111;
				8'b1000111: c <= 9'b110001111;
				8'b1011111: c <= 9'b11011001;
				8'b1110100: c <= 9'b11100011;
				8'b101101: c <= 9'b10101100;
				8'b1010011: c <= 9'b1010110;
				8'b1100001: c <= 9'b1001;
				8'b110101: c <= 9'b110010011;
				8'b1000100: c <= 9'b110001110;
				8'b1010001: c <= 9'b10110100;
				8'b1010100: c <= 9'b100011101;
				8'b1100110: c <= 9'b101000;
				8'b101010: c <= 9'b101000100;
				8'b1011110: c <= 9'b11011001;
				8'b1100111: c <= 9'b11000110;
				8'b1011010: c <= 9'b11111101;
				8'b1000010: c <= 9'b10011;
				8'b111101: c <= 9'b111010110;
				8'b110000: c <= 9'b111111011;
				8'b111110: c <= 9'b10010111;
				8'b1100010: c <= 9'b1001010;
				8'b1110000: c <= 9'b1000111;
				8'b1101001: c <= 9'b110001;
				8'b1110011: c <= 9'b11010111;
				8'b1001100: c <= 9'b101101010;
				8'b100001: c <= 9'b100111010;
				8'b1000110: c <= 9'b101001001;
				8'b1110010: c <= 9'b111001;
				8'b1010000: c <= 9'b110011101;
				8'b1111010: c <= 9'b1000111;
				8'b1010101: c <= 9'b101011011;
				8'b111011: c <= 9'b11101101;
				8'b1001101: c <= 9'b111100010;
				8'b111111: c <= 9'b11111;
				8'b1101110: c <= 9'b1010001;
				8'b1111011: c <= 9'b101101001;
				8'b1001011: c <= 9'b1010110;
				8'b1101111: c <= 9'b1111111;
				8'b1101000: c <= 9'b101100;
				8'b101100: c <= 9'b1010010;
				8'b100100: c <= 9'b11011101;
				8'b1111000: c <= 9'b110111100;
				8'b1000101: c <= 9'b10101;
				8'b1011001: c <= 9'b111100111;
				8'b110100: c <= 9'b1000101;
				8'b1111001: c <= 9'b101111000;
				8'b1110001: c <= 9'b100010000;
				8'b1001111: c <= 9'b1111001;
				8'b1100101: c <= 9'b101001001;
				8'b1111110: c <= 9'b1100101;
				8'b1111100: c <= 9'b111011010;
				8'b1010110: c <= 9'b101101010;
				8'b110010: c <= 9'b111011;
				8'b1101101: c <= 9'b101101011;
				8'b100011: c <= 9'b111111010;
				8'b1110101: c <= 9'b110001101;
				8'b1111101: c <= 9'b101011;
				8'b101001: c <= 9'b100111001;
				8'b1010010: c <= 9'b100101001;
				8'b1011000: c <= 9'b11011011;
				8'b101110: c <= 9'b11101100;
				8'b1000001: c <= 9'b10101101;
				default: c <= 9'b0;
			endcase
			9'b10001100 : case(di)
				8'b1000011: c <= 9'b111001010;
				8'b101000: c <= 9'b110000011;
				8'b111010: c <= 9'b110000001;
				8'b110110: c <= 9'b100101001;
				8'b1100100: c <= 9'b11011110;
				8'b1000000: c <= 9'b1111101;
				8'b1110110: c <= 9'b111111011;
				8'b100101: c <= 9'b101110101;
				8'b101111: c <= 9'b100100010;
				8'b100110: c <= 9'b11;
				8'b1100011: c <= 9'b100000011;
				8'b1001000: c <= 9'b111111101;
				8'b111000: c <= 9'b1001010;
				8'b110001: c <= 9'b101100000;
				8'b1010111: c <= 9'b111001010;
				8'b1001110: c <= 9'b11100000;
				8'b1101010: c <= 9'b111101110;
				8'b1001001: c <= 9'b100010011;
				8'b1100000: c <= 9'b11001100;
				8'b110111: c <= 9'b110110011;
				8'b1011101: c <= 9'b100110010;
				8'b1011011: c <= 9'b10100111;
				8'b111001: c <= 9'b101010011;
				8'b1001010: c <= 9'b110100010;
				8'b110011: c <= 9'b1101;
				8'b1101100: c <= 9'b100001;
				8'b1110111: c <= 9'b11111100;
				8'b101011: c <= 9'b1010010;
				8'b1101011: c <= 9'b110110;
				8'b111100: c <= 9'b1100000;
				8'b1000111: c <= 9'b11011010;
				8'b1011111: c <= 9'b101010010;
				8'b1110100: c <= 9'b100101101;
				8'b101101: c <= 9'b100110;
				8'b1010011: c <= 9'b111100011;
				8'b1100001: c <= 9'b100101001;
				8'b110101: c <= 9'b100000111;
				8'b1000100: c <= 9'b111101000;
				8'b1010001: c <= 9'b111111010;
				8'b1010100: c <= 9'b110100100;
				8'b1100110: c <= 9'b110011011;
				8'b101010: c <= 9'b100101100;
				8'b1011110: c <= 9'b1010011;
				8'b1100111: c <= 9'b100001100;
				8'b1011010: c <= 9'b1101110;
				8'b1000010: c <= 9'b101100100;
				8'b111101: c <= 9'b1111110;
				8'b110000: c <= 9'b11001111;
				8'b111110: c <= 9'b10110111;
				8'b1100010: c <= 9'b11111010;
				8'b1110000: c <= 9'b111000100;
				8'b1101001: c <= 9'b10010100;
				8'b1110011: c <= 9'b11000100;
				8'b1001100: c <= 9'b10101100;
				8'b100001: c <= 9'b10000110;
				8'b1000110: c <= 9'b110001010;
				8'b1110010: c <= 9'b100010011;
				8'b1010000: c <= 9'b10001101;
				8'b1111010: c <= 9'b111101101;
				8'b1010101: c <= 9'b101000011;
				8'b111011: c <= 9'b111000111;
				8'b1001101: c <= 9'b110011101;
				8'b111111: c <= 9'b10011;
				8'b1101110: c <= 9'b10101001;
				8'b1111011: c <= 9'b101101100;
				8'b1001011: c <= 9'b1001000;
				8'b1101111: c <= 9'b11010;
				8'b1101000: c <= 9'b1000010;
				8'b101100: c <= 9'b100101101;
				8'b100100: c <= 9'b101011000;
				8'b1111000: c <= 9'b101;
				8'b1000101: c <= 9'b1111011;
				8'b1011001: c <= 9'b111001110;
				8'b110100: c <= 9'b1001001;
				8'b1111001: c <= 9'b111001010;
				8'b1110001: c <= 9'b111001000;
				8'b1001111: c <= 9'b101111010;
				8'b1100101: c <= 9'b10001010;
				8'b1111110: c <= 9'b101101101;
				8'b1111100: c <= 9'b100111100;
				8'b1010110: c <= 9'b101110010;
				8'b110010: c <= 9'b1000001;
				8'b1101101: c <= 9'b100011100;
				8'b100011: c <= 9'b100101101;
				8'b1110101: c <= 9'b1010111;
				8'b1111101: c <= 9'b111011100;
				8'b101001: c <= 9'b1011010;
				8'b1010010: c <= 9'b100000010;
				8'b1011000: c <= 9'b100111001;
				8'b101110: c <= 9'b101111111;
				8'b1000001: c <= 9'b111110001;
				default: c <= 9'b0;
			endcase
			9'b11100000 : case(di)
				8'b1000011: c <= 9'b10111100;
				8'b101000: c <= 9'b1101001;
				8'b111010: c <= 9'b111010;
				8'b110110: c <= 9'b110010100;
				8'b1100100: c <= 9'b110100;
				8'b1000000: c <= 9'b111000110;
				8'b1110110: c <= 9'b111001000;
				8'b100101: c <= 9'b11110001;
				8'b101111: c <= 9'b111001101;
				8'b100110: c <= 9'b11111100;
				8'b1100011: c <= 9'b1101000;
				8'b1001000: c <= 9'b110011110;
				8'b111000: c <= 9'b100101;
				8'b110001: c <= 9'b10001110;
				8'b1010111: c <= 9'b1101100;
				8'b1001110: c <= 9'b110101101;
				8'b1101010: c <= 9'b1100100;
				8'b1001001: c <= 9'b1000000;
				8'b1100000: c <= 9'b100001110;
				8'b110111: c <= 9'b100000001;
				8'b1011101: c <= 9'b10110110;
				8'b1011011: c <= 9'b1101001;
				8'b111001: c <= 9'b110111110;
				8'b1001010: c <= 9'b110000000;
				8'b110011: c <= 9'b110011011;
				8'b1101100: c <= 9'b100111001;
				8'b1110111: c <= 9'b111110000;
				8'b101011: c <= 9'b111100100;
				8'b1101011: c <= 9'b110011001;
				8'b111100: c <= 9'b110110011;
				8'b1000111: c <= 9'b100000100;
				8'b1011111: c <= 9'b110101001;
				8'b1110100: c <= 9'b110101011;
				8'b101101: c <= 9'b1;
				8'b1010011: c <= 9'b111101000;
				8'b1100001: c <= 9'b100110;
				8'b110101: c <= 9'b10100;
				8'b1000100: c <= 9'b10100100;
				8'b1010001: c <= 9'b110110;
				8'b1010100: c <= 9'b10100;
				8'b1100110: c <= 9'b1100101;
				8'b101010: c <= 9'b1100100;
				8'b1011110: c <= 9'b100000000;
				8'b1100111: c <= 9'b101010101;
				8'b1011010: c <= 9'b110001100;
				8'b1000010: c <= 9'b10010001;
				8'b111101: c <= 9'b101101000;
				8'b110000: c <= 9'b10000010;
				8'b111110: c <= 9'b110100010;
				8'b1100010: c <= 9'b10011010;
				8'b1110000: c <= 9'b1011011;
				8'b1101001: c <= 9'b10010;
				8'b1110011: c <= 9'b110100100;
				8'b1001100: c <= 9'b101010111;
				8'b100001: c <= 9'b10000010;
				8'b1000110: c <= 9'b110111000;
				8'b1110010: c <= 9'b101100000;
				8'b1010000: c <= 9'b101100001;
				8'b1111010: c <= 9'b11010011;
				8'b1010101: c <= 9'b111101110;
				8'b111011: c <= 9'b100100010;
				8'b1001101: c <= 9'b1101010;
				8'b111111: c <= 9'b10011010;
				8'b1101110: c <= 9'b1101000;
				8'b1111011: c <= 9'b111111010;
				8'b1001011: c <= 9'b111111101;
				8'b1101111: c <= 9'b101100;
				8'b1101000: c <= 9'b10110110;
				8'b101100: c <= 9'b101000001;
				8'b100100: c <= 9'b111;
				8'b1111000: c <= 9'b101001000;
				8'b1000101: c <= 9'b10001110;
				8'b1011001: c <= 9'b100000011;
				8'b110100: c <= 9'b100011101;
				8'b1111001: c <= 9'b110011000;
				8'b1110001: c <= 9'b11001001;
				8'b1001111: c <= 9'b110010100;
				8'b1100101: c <= 9'b111111101;
				8'b1111110: c <= 9'b101110100;
				8'b1111100: c <= 9'b100011101;
				8'b1010110: c <= 9'b11111101;
				8'b110010: c <= 9'b100111;
				8'b1101101: c <= 9'b100100010;
				8'b100011: c <= 9'b101101011;
				8'b1110101: c <= 9'b10000010;
				8'b1111101: c <= 9'b10101010;
				8'b101001: c <= 9'b11110101;
				8'b1010010: c <= 9'b101000100;
				8'b1011000: c <= 9'b101000101;
				8'b101110: c <= 9'b11100011;
				8'b1000001: c <= 9'b111110000;
				default: c <= 9'b0;
			endcase
			9'b100101100 : case(di)
				8'b1000011: c <= 9'b11011110;
				8'b101000: c <= 9'b100111001;
				8'b111010: c <= 9'b10001011;
				8'b110110: c <= 9'b11100;
				8'b1100100: c <= 9'b111101010;
				8'b1000000: c <= 9'b111101000;
				8'b1110110: c <= 9'b111001110;
				8'b100101: c <= 9'b10100110;
				8'b101111: c <= 9'b110100;
				8'b100110: c <= 9'b111001110;
				8'b1100011: c <= 9'b10010100;
				8'b1001000: c <= 9'b101110100;
				8'b111000: c <= 9'b10000101;
				8'b110001: c <= 9'b10110111;
				8'b1010111: c <= 9'b111000111;
				8'b1001110: c <= 9'b101110110;
				8'b1101010: c <= 9'b101001010;
				8'b1001001: c <= 9'b101111111;
				8'b1100000: c <= 9'b100001;
				8'b110111: c <= 9'b110001100;
				8'b1011101: c <= 9'b100010010;
				8'b1011011: c <= 9'b100100;
				8'b111001: c <= 9'b111111111;
				8'b1001010: c <= 9'b1100010;
				8'b110011: c <= 9'b100101101;
				8'b1101100: c <= 9'b110110010;
				8'b1110111: c <= 9'b11010100;
				8'b101011: c <= 9'b110000010;
				8'b1101011: c <= 9'b110110000;
				8'b111100: c <= 9'b101101011;
				8'b1000111: c <= 9'b1011100;
				8'b1011111: c <= 9'b101001110;
				8'b1110100: c <= 9'b1110000;
				8'b101101: c <= 9'b101000011;
				8'b1010011: c <= 9'b100111011;
				8'b1100001: c <= 9'b101100110;
				8'b110101: c <= 9'b111000101;
				8'b1000100: c <= 9'b110010100;
				8'b1010001: c <= 9'b101011111;
				8'b1010100: c <= 9'b111010111;
				8'b1100110: c <= 9'b10110101;
				8'b101010: c <= 9'b111100101;
				8'b1011110: c <= 9'b10010111;
				8'b1100111: c <= 9'b11110010;
				8'b1011010: c <= 9'b100000100;
				8'b1000010: c <= 9'b1111001;
				8'b111101: c <= 9'b1010000;
				8'b110000: c <= 9'b101110011;
				8'b111110: c <= 9'b111001100;
				8'b1100010: c <= 9'b11;
				8'b1110000: c <= 9'b110101010;
				8'b1101001: c <= 9'b110101010;
				8'b1110011: c <= 9'b10010001;
				8'b1001100: c <= 9'b1001;
				8'b100001: c <= 9'b111000100;
				8'b1000110: c <= 9'b101011000;
				8'b1110010: c <= 9'b11001010;
				8'b1010000: c <= 9'b11001100;
				8'b1111010: c <= 9'b101100000;
				8'b1010101: c <= 9'b10111100;
				8'b111011: c <= 9'b100101100;
				8'b1001101: c <= 9'b110110111;
				8'b111111: c <= 9'b110110000;
				8'b1101110: c <= 9'b11101;
				8'b1111011: c <= 9'b111101010;
				8'b1001011: c <= 9'b10110010;
				8'b1101111: c <= 9'b111001001;
				8'b1101000: c <= 9'b110111000;
				8'b101100: c <= 9'b1110011;
				8'b100100: c <= 9'b100011010;
				8'b1111000: c <= 9'b100100011;
				8'b1000101: c <= 9'b100000010;
				8'b1011001: c <= 9'b100010010;
				8'b110100: c <= 9'b10101010;
				8'b1111001: c <= 9'b11010001;
				8'b1110001: c <= 9'b110111011;
				8'b1001111: c <= 9'b1111111;
				8'b1100101: c <= 9'b111111011;
				8'b1111110: c <= 9'b1000100;
				8'b1111100: c <= 9'b11010010;
				8'b1010110: c <= 9'b1101000;
				8'b110010: c <= 9'b100100001;
				8'b1101101: c <= 9'b11011011;
				8'b100011: c <= 9'b101010;
				8'b1110101: c <= 9'b110111100;
				8'b1111101: c <= 9'b11010010;
				8'b101001: c <= 9'b10010000;
				8'b1010010: c <= 9'b101011111;
				8'b1011000: c <= 9'b100111111;
				8'b101110: c <= 9'b10000010;
				8'b1000001: c <= 9'b101101011;
				default: c <= 9'b0;
			endcase
			9'b10110111 : case(di)
				8'b1000011: c <= 9'b111000000;
				8'b101000: c <= 9'b100000111;
				8'b111010: c <= 9'b1100101;
				8'b110110: c <= 9'b111111011;
				8'b1100100: c <= 9'b1000110;
				8'b1000000: c <= 9'b111001111;
				8'b1110110: c <= 9'b11010001;
				8'b100101: c <= 9'b111010100;
				8'b101111: c <= 9'b110000001;
				8'b100110: c <= 9'b111100110;
				8'b1100011: c <= 9'b10001110;
				8'b1001000: c <= 9'b101110100;
				8'b111000: c <= 9'b11100001;
				8'b110001: c <= 9'b101110;
				8'b1010111: c <= 9'b10100011;
				8'b1001110: c <= 9'b10011100;
				8'b1101010: c <= 9'b11001101;
				8'b1001001: c <= 9'b10101;
				8'b1100000: c <= 9'b101001110;
				8'b110111: c <= 9'b11111101;
				8'b1011101: c <= 9'b101010101;
				8'b1011011: c <= 9'b100000101;
				8'b111001: c <= 9'b111011;
				8'b1001010: c <= 9'b11000011;
				8'b110011: c <= 9'b1110;
				8'b1101100: c <= 9'b100011011;
				8'b1110111: c <= 9'b1101000;
				8'b101011: c <= 9'b101101001;
				8'b1101011: c <= 9'b10011010;
				8'b111100: c <= 9'b10110;
				8'b1000111: c <= 9'b111100001;
				8'b1011111: c <= 9'b111010000;
				8'b1110100: c <= 9'b11001111;
				8'b101101: c <= 9'b111110011;
				8'b1010011: c <= 9'b11000111;
				8'b1100001: c <= 9'b100001;
				8'b110101: c <= 9'b100111001;
				8'b1000100: c <= 9'b111100101;
				8'b1010001: c <= 9'b1110100;
				8'b1010100: c <= 9'b111101111;
				8'b1100110: c <= 9'b111001001;
				8'b101010: c <= 9'b111001110;
				8'b1011110: c <= 9'b1100100;
				8'b1100111: c <= 9'b1001110;
				8'b1011010: c <= 9'b110111110;
				8'b1000010: c <= 9'b100010;
				8'b111101: c <= 9'b100100011;
				8'b110000: c <= 9'b101110100;
				8'b111110: c <= 9'b100010110;
				8'b1100010: c <= 9'b11100011;
				8'b1110000: c <= 9'b100111111;
				8'b1101001: c <= 9'b11010001;
				8'b1110011: c <= 9'b1110100;
				8'b1001100: c <= 9'b101011001;
				8'b100001: c <= 9'b101011111;
				8'b1000110: c <= 9'b10010111;
				8'b1110010: c <= 9'b10100110;
				8'b1010000: c <= 9'b1111101;
				8'b1111010: c <= 9'b11101101;
				8'b1010101: c <= 9'b100110011;
				8'b111011: c <= 9'b100010;
				8'b1001101: c <= 9'b110001111;
				8'b111111: c <= 9'b110100000;
				8'b1101110: c <= 9'b101101101;
				8'b1111011: c <= 9'b110100100;
				8'b1001011: c <= 9'b1001010;
				8'b1101111: c <= 9'b110110100;
				8'b1101000: c <= 9'b1010110;
				8'b101100: c <= 9'b101001010;
				8'b100100: c <= 9'b1101110;
				8'b1111000: c <= 9'b11010010;
				8'b1000101: c <= 9'b101010100;
				8'b1011001: c <= 9'b101100101;
				8'b110100: c <= 9'b110010010;
				8'b1111001: c <= 9'b10111101;
				8'b1110001: c <= 9'b110101001;
				8'b1001111: c <= 9'b110111000;
				8'b1100101: c <= 9'b110010111;
				8'b1111110: c <= 9'b100100;
				8'b1111100: c <= 9'b101011101;
				8'b1010110: c <= 9'b111100000;
				8'b110010: c <= 9'b1111110;
				8'b1101101: c <= 9'b101001011;
				8'b100011: c <= 9'b1000100;
				8'b1110101: c <= 9'b111101111;
				8'b1111101: c <= 9'b10110;
				8'b101001: c <= 9'b100001100;
				8'b1010010: c <= 9'b10111000;
				8'b1011000: c <= 9'b11110000;
				8'b101110: c <= 9'b1000;
				8'b1000001: c <= 9'b100001011;
				default: c <= 9'b0;
			endcase
			9'b11110011 : case(di)
				8'b1000011: c <= 9'b100;
				8'b101000: c <= 9'b111000101;
				8'b111010: c <= 9'b11101101;
				8'b110110: c <= 9'b1011011;
				8'b1100100: c <= 9'b101100110;
				8'b1000000: c <= 9'b110011011;
				8'b1110110: c <= 9'b101001011;
				8'b100101: c <= 9'b111101100;
				8'b101111: c <= 9'b11001;
				8'b100110: c <= 9'b100110100;
				8'b1100011: c <= 9'b10001100;
				8'b1001000: c <= 9'b110001001;
				8'b111000: c <= 9'b110001110;
				8'b110001: c <= 9'b10110100;
				8'b1010111: c <= 9'b1110001;
				8'b1001110: c <= 9'b101010010;
				8'b1101010: c <= 9'b10001000;
				8'b1001001: c <= 9'b110100010;
				8'b1100000: c <= 9'b10011011;
				8'b110111: c <= 9'b11010011;
				8'b1011101: c <= 9'b10100100;
				8'b1011011: c <= 9'b100111101;
				8'b111001: c <= 9'b111001110;
				8'b1001010: c <= 9'b100111000;
				8'b110011: c <= 9'b10101001;
				8'b1101100: c <= 9'b100110101;
				8'b1110111: c <= 9'b11000000;
				8'b101011: c <= 9'b111110001;
				8'b1101011: c <= 9'b11100100;
				8'b111100: c <= 9'b1010011;
				8'b1000111: c <= 9'b111010001;
				8'b1011111: c <= 9'b111110001;
				8'b1110100: c <= 9'b111000110;
				8'b101101: c <= 9'b111011111;
				8'b1010011: c <= 9'b10010111;
				8'b1100001: c <= 9'b101111110;
				8'b110101: c <= 9'b110100011;
				8'b1000100: c <= 9'b100111100;
				8'b1010001: c <= 9'b100011100;
				8'b1010100: c <= 9'b100010100;
				8'b1100110: c <= 9'b1110010;
				8'b101010: c <= 9'b100001011;
				8'b1011110: c <= 9'b10001100;
				8'b1100111: c <= 9'b100111101;
				8'b1011010: c <= 9'b10000101;
				8'b1000010: c <= 9'b1001100;
				8'b111101: c <= 9'b111101110;
				8'b110000: c <= 9'b111001000;
				8'b111110: c <= 9'b100000100;
				8'b1100010: c <= 9'b1001101;
				8'b1110000: c <= 9'b100011111;
				8'b1101001: c <= 9'b100100000;
				8'b1110011: c <= 9'b101111001;
				8'b1001100: c <= 9'b111101101;
				8'b100001: c <= 9'b11000110;
				8'b1000110: c <= 9'b110101101;
				8'b1110010: c <= 9'b110010011;
				8'b1010000: c <= 9'b111000100;
				8'b1111010: c <= 9'b111111101;
				8'b1010101: c <= 9'b10101100;
				8'b111011: c <= 9'b111111001;
				8'b1001101: c <= 9'b110000001;
				8'b111111: c <= 9'b1101001;
				8'b1101110: c <= 9'b110110;
				8'b1111011: c <= 9'b1011;
				8'b1001011: c <= 9'b101000;
				8'b1101111: c <= 9'b100011011;
				8'b1101000: c <= 9'b11111110;
				8'b101100: c <= 9'b10000010;
				8'b100100: c <= 9'b11010111;
				8'b1111000: c <= 9'b110000010;
				8'b1000101: c <= 9'b11010;
				8'b1011001: c <= 9'b101010001;
				8'b110100: c <= 9'b100010;
				8'b1111001: c <= 9'b1011;
				8'b1110001: c <= 9'b10101100;
				8'b1001111: c <= 9'b110000101;
				8'b1100101: c <= 9'b110000111;
				8'b1111110: c <= 9'b101001001;
				8'b1111100: c <= 9'b100000010;
				8'b1010110: c <= 9'b100010011;
				8'b110010: c <= 9'b100011001;
				8'b1101101: c <= 9'b100000111;
				8'b100011: c <= 9'b110110100;
				8'b1110101: c <= 9'b11000;
				8'b1111101: c <= 9'b100111110;
				8'b101001: c <= 9'b1010010;
				8'b1010010: c <= 9'b110011110;
				8'b1011000: c <= 9'b101001001;
				8'b101110: c <= 9'b100000000;
				8'b1000001: c <= 9'b101001001;
				default: c <= 9'b0;
			endcase
			9'b100000000 : case(di)
				8'b1000011: c <= 9'b111100011;
				8'b101000: c <= 9'b11100;
				8'b111010: c <= 9'b11101101;
				8'b110110: c <= 9'b1010111;
				8'b1100100: c <= 9'b110110010;
				8'b1000000: c <= 9'b10111110;
				8'b1110110: c <= 9'b101110010;
				8'b100101: c <= 9'b101001111;
				8'b101111: c <= 9'b100011100;
				8'b100110: c <= 9'b1000100;
				8'b1100011: c <= 9'b100001011;
				8'b1001000: c <= 9'b110111001;
				8'b111000: c <= 9'b111000111;
				8'b110001: c <= 9'b110111110;
				8'b1010111: c <= 9'b1010110;
				8'b1001110: c <= 9'b100100111;
				8'b1101010: c <= 9'b101100;
				8'b1001001: c <= 9'b110010110;
				8'b1100000: c <= 9'b101000110;
				8'b110111: c <= 9'b100010101;
				8'b1011101: c <= 9'b110100101;
				8'b1011011: c <= 9'b101111000;
				8'b111001: c <= 9'b110111100;
				8'b1001010: c <= 9'b101011001;
				8'b110011: c <= 9'b10000011;
				8'b1101100: c <= 9'b11111001;
				8'b1110111: c <= 9'b110011111;
				8'b101011: c <= 9'b11010000;
				8'b1101011: c <= 9'b101100001;
				8'b111100: c <= 9'b110001011;
				8'b1000111: c <= 9'b111110110;
				8'b1011111: c <= 9'b100100;
				8'b1110100: c <= 9'b11001111;
				8'b101101: c <= 9'b111101101;
				8'b1010011: c <= 9'b111111001;
				8'b1100001: c <= 9'b10001110;
				8'b110101: c <= 9'b11000;
				8'b1000100: c <= 9'b11111010;
				8'b1010001: c <= 9'b110011011;
				8'b1010100: c <= 9'b101011000;
				8'b1100110: c <= 9'b101010;
				8'b101010: c <= 9'b110110011;
				8'b1011110: c <= 9'b101100011;
				8'b1100111: c <= 9'b10;
				8'b1011010: c <= 9'b1000011;
				8'b1000010: c <= 9'b101001110;
				8'b111101: c <= 9'b1000000;
				8'b110000: c <= 9'b10111000;
				8'b111110: c <= 9'b101110001;
				8'b1100010: c <= 9'b100000101;
				8'b1110000: c <= 9'b1001110;
				8'b1101001: c <= 9'b100011011;
				8'b1110011: c <= 9'b1101110;
				8'b1001100: c <= 9'b111111;
				8'b100001: c <= 9'b11100100;
				8'b1000110: c <= 9'b100011101;
				8'b1110010: c <= 9'b110001111;
				8'b1010000: c <= 9'b10000011;
				8'b1111010: c <= 9'b100010001;
				8'b1010101: c <= 9'b101011011;
				8'b111011: c <= 9'b110011111;
				8'b1001101: c <= 9'b1010010;
				8'b111111: c <= 9'b10;
				8'b1101110: c <= 9'b111101;
				8'b1111011: c <= 9'b111100101;
				8'b1001011: c <= 9'b100011100;
				8'b1101111: c <= 9'b101100001;
				8'b1101000: c <= 9'b110010011;
				8'b101100: c <= 9'b11111;
				8'b100100: c <= 9'b10001110;
				8'b1111000: c <= 9'b100100001;
				8'b1000101: c <= 9'b10100111;
				8'b1011001: c <= 9'b111011001;
				8'b110100: c <= 9'b1110;
				8'b1111001: c <= 9'b110011101;
				8'b1110001: c <= 9'b11100000;
				8'b1001111: c <= 9'b1100100;
				8'b1100101: c <= 9'b1100101;
				8'b1111110: c <= 9'b110000110;
				8'b1111100: c <= 9'b100000110;
				8'b1010110: c <= 9'b100111100;
				8'b110010: c <= 9'b110011011;
				8'b1101101: c <= 9'b110010001;
				8'b100011: c <= 9'b100000101;
				8'b1110101: c <= 9'b10101001;
				8'b1111101: c <= 9'b11110000;
				8'b101001: c <= 9'b110010111;
				8'b1010010: c <= 9'b1100000;
				8'b1011000: c <= 9'b110001;
				8'b101110: c <= 9'b111001110;
				8'b1000001: c <= 9'b1110;
				default: c <= 9'b0;
			endcase
			9'b11111000 : case(di)
				8'b1000011: c <= 9'b101101011;
				8'b101000: c <= 9'b100101010;
				8'b111010: c <= 9'b101111010;
				8'b110110: c <= 9'b101010010;
				8'b1100100: c <= 9'b101111110;
				8'b1000000: c <= 9'b1101000;
				8'b1110110: c <= 9'b100111110;
				8'b100101: c <= 9'b111011010;
				8'b101111: c <= 9'b101100100;
				8'b100110: c <= 9'b11001111;
				8'b1100011: c <= 9'b10001101;
				8'b1001000: c <= 9'b10101111;
				8'b111000: c <= 9'b1111110;
				8'b110001: c <= 9'b111100110;
				8'b1010111: c <= 9'b10000;
				8'b1001110: c <= 9'b101011010;
				8'b1101010: c <= 9'b1011100;
				8'b1001001: c <= 9'b111001;
				8'b1100000: c <= 9'b111001010;
				8'b110111: c <= 9'b111110110;
				8'b1011101: c <= 9'b11111;
				8'b1011011: c <= 9'b1001001;
				8'b111001: c <= 9'b100110101;
				8'b1001010: c <= 9'b1111100;
				8'b110011: c <= 9'b110101011;
				8'b1101100: c <= 9'b101001100;
				8'b1110111: c <= 9'b11010001;
				8'b101011: c <= 9'b101011001;
				8'b1101011: c <= 9'b10111110;
				8'b111100: c <= 9'b111111011;
				8'b1000111: c <= 9'b101001001;
				8'b1011111: c <= 9'b111101010;
				8'b1110100: c <= 9'b10101100;
				8'b101101: c <= 9'b11001100;
				8'b1010011: c <= 9'b111011110;
				8'b1100001: c <= 9'b1000101;
				8'b110101: c <= 9'b1101000;
				8'b1000100: c <= 9'b100101000;
				8'b1010001: c <= 9'b101111001;
				8'b1010100: c <= 9'b10;
				8'b1100110: c <= 9'b111101100;
				8'b101010: c <= 9'b1111100;
				8'b1011110: c <= 9'b1110000;
				8'b1100111: c <= 9'b111001010;
				8'b1011010: c <= 9'b11100110;
				8'b1000010: c <= 9'b101100001;
				8'b111101: c <= 9'b11001010;
				8'b110000: c <= 9'b10100100;
				8'b111110: c <= 9'b10100000;
				8'b1100010: c <= 9'b1100;
				8'b1110000: c <= 9'b100001111;
				8'b1101001: c <= 9'b101000;
				8'b1110011: c <= 9'b10101;
				8'b1001100: c <= 9'b110000000;
				8'b100001: c <= 9'b10011;
				8'b1000110: c <= 9'b11001;
				8'b1110010: c <= 9'b11111100;
				8'b1010000: c <= 9'b110101001;
				8'b1111010: c <= 9'b10111110;
				8'b1010101: c <= 9'b10111;
				8'b111011: c <= 9'b101100101;
				8'b1001101: c <= 9'b10001011;
				8'b111111: c <= 9'b11000000;
				8'b1101110: c <= 9'b110101;
				8'b1111011: c <= 9'b100101010;
				8'b1001011: c <= 9'b1011;
				8'b1101111: c <= 9'b1010010;
				8'b1101000: c <= 9'b11100011;
				8'b101100: c <= 9'b101011111;
				8'b100100: c <= 9'b10110;
				8'b1111000: c <= 9'b10100011;
				8'b1000101: c <= 9'b100101110;
				8'b1011001: c <= 9'b110010111;
				8'b110100: c <= 9'b101000100;
				8'b1111001: c <= 9'b100001111;
				8'b1110001: c <= 9'b11000100;
				8'b1001111: c <= 9'b10111000;
				8'b1100101: c <= 9'b10111111;
				8'b1111110: c <= 9'b111000011;
				8'b1111100: c <= 9'b101101010;
				8'b1010110: c <= 9'b101101000;
				8'b110010: c <= 9'b11110100;
				8'b1101101: c <= 9'b101101010;
				8'b100011: c <= 9'b110000010;
				8'b1110101: c <= 9'b11101011;
				8'b1111101: c <= 9'b111100;
				8'b101001: c <= 9'b11110011;
				8'b1010010: c <= 9'b110010101;
				8'b1011000: c <= 9'b111011010;
				8'b101110: c <= 9'b1010111;
				8'b1000001: c <= 9'b1111;
				default: c <= 9'b0;
			endcase
			9'b100100010 : case(di)
				8'b1000011: c <= 9'b11001111;
				8'b101000: c <= 9'b111111101;
				8'b111010: c <= 9'b10111001;
				8'b110110: c <= 9'b100010;
				8'b1100100: c <= 9'b11101000;
				8'b1000000: c <= 9'b101100110;
				8'b1110110: c <= 9'b100101011;
				8'b100101: c <= 9'b10101101;
				8'b101111: c <= 9'b1101010;
				8'b100110: c <= 9'b11101001;
				8'b1100011: c <= 9'b101111000;
				8'b1001000: c <= 9'b100101111;
				8'b111000: c <= 9'b10100100;
				8'b110001: c <= 9'b11100101;
				8'b1010111: c <= 9'b10110010;
				8'b1001110: c <= 9'b111010001;
				8'b1101010: c <= 9'b10101011;
				8'b1001001: c <= 9'b100111010;
				8'b1100000: c <= 9'b101110100;
				8'b110111: c <= 9'b101001111;
				8'b1011101: c <= 9'b111101110;
				8'b1011011: c <= 9'b111001110;
				8'b111001: c <= 9'b10101111;
				8'b1001010: c <= 9'b111111001;
				8'b110011: c <= 9'b111000011;
				8'b1101100: c <= 9'b100111001;
				8'b1110111: c <= 9'b101100;
				8'b101011: c <= 9'b101101;
				8'b1101011: c <= 9'b111111101;
				8'b111100: c <= 9'b11101;
				8'b1000111: c <= 9'b1101100;
				8'b1011111: c <= 9'b1110000;
				8'b1110100: c <= 9'b100110;
				8'b101101: c <= 9'b101101100;
				8'b1010011: c <= 9'b101011001;
				8'b1100001: c <= 9'b11000011;
				8'b110101: c <= 9'b1000101;
				8'b1000100: c <= 9'b1101111;
				8'b1010001: c <= 9'b10000111;
				8'b1010100: c <= 9'b101101010;
				8'b1100110: c <= 9'b100110111;
				8'b101010: c <= 9'b111110110;
				8'b1011110: c <= 9'b100000100;
				8'b1100111: c <= 9'b101011101;
				8'b1011010: c <= 9'b110000000;
				8'b1000010: c <= 9'b10111001;
				8'b111101: c <= 9'b100101110;
				8'b110000: c <= 9'b101110100;
				8'b111110: c <= 9'b11111001;
				8'b1100010: c <= 9'b1100000;
				8'b1110000: c <= 9'b110001111;
				8'b1101001: c <= 9'b110010100;
				8'b1110011: c <= 9'b110110110;
				8'b1001100: c <= 9'b101110011;
				8'b100001: c <= 9'b111011001;
				8'b1000110: c <= 9'b111001100;
				8'b1110010: c <= 9'b1101001;
				8'b1010000: c <= 9'b101010000;
				8'b1111010: c <= 9'b110100001;
				8'b1010101: c <= 9'b100111;
				8'b111011: c <= 9'b11001111;
				8'b1001101: c <= 9'b11001011;
				8'b111111: c <= 9'b11101100;
				8'b1101110: c <= 9'b100;
				8'b1111011: c <= 9'b11000;
				8'b1001011: c <= 9'b10101011;
				8'b1101111: c <= 9'b1100001;
				8'b1101000: c <= 9'b100001011;
				8'b101100: c <= 9'b11011110;
				8'b100100: c <= 9'b111001111;
				8'b1111000: c <= 9'b1011001;
				8'b1000101: c <= 9'b110100100;
				8'b1011001: c <= 9'b100001110;
				8'b110100: c <= 9'b111100011;
				8'b1111001: c <= 9'b110000000;
				8'b1110001: c <= 9'b1100110;
				8'b1001111: c <= 9'b100011100;
				8'b1100101: c <= 9'b110100001;
				8'b1111110: c <= 9'b100110011;
				8'b1111100: c <= 9'b101000101;
				8'b1010110: c <= 9'b110010001;
				8'b110010: c <= 9'b100000010;
				8'b1101101: c <= 9'b110111001;
				8'b100011: c <= 9'b11001101;
				8'b1110101: c <= 9'b10101;
				8'b1111101: c <= 9'b111001;
				8'b101001: c <= 9'b10110110;
				8'b1010010: c <= 9'b100110101;
				8'b1011000: c <= 9'b101110111;
				8'b101110: c <= 9'b1011110;
				8'b1000001: c <= 9'b10001110;
				default: c <= 9'b0;
			endcase
			9'b11010100 : case(di)
				8'b1000011: c <= 9'b110001011;
				8'b101000: c <= 9'b101100111;
				8'b111010: c <= 9'b101011011;
				8'b110110: c <= 9'b10010;
				8'b1100100: c <= 9'b111011010;
				8'b1000000: c <= 9'b110010101;
				8'b1110110: c <= 9'b110100011;
				8'b100101: c <= 9'b100101111;
				8'b101111: c <= 9'b1100100;
				8'b100110: c <= 9'b101001001;
				8'b1100011: c <= 9'b100010011;
				8'b1001000: c <= 9'b111100011;
				8'b111000: c <= 9'b10101000;
				8'b110001: c <= 9'b100111011;
				8'b1010111: c <= 9'b110001100;
				8'b1001110: c <= 9'b11010001;
				8'b1101010: c <= 9'b1101111;
				8'b1001001: c <= 9'b11100;
				8'b1100000: c <= 9'b1101110;
				8'b110111: c <= 9'b1001001;
				8'b1011101: c <= 9'b110011000;
				8'b1011011: c <= 9'b110110;
				8'b111001: c <= 9'b110101011;
				8'b1001010: c <= 9'b110100001;
				8'b110011: c <= 9'b1111111;
				8'b1101100: c <= 9'b110001001;
				8'b1110111: c <= 9'b1110000;
				8'b101011: c <= 9'b110110101;
				8'b1101011: c <= 9'b10101100;
				8'b111100: c <= 9'b11011011;
				8'b1000111: c <= 9'b111011110;
				8'b1011111: c <= 9'b1101010;
				8'b1110100: c <= 9'b101110000;
				8'b101101: c <= 9'b100110010;
				8'b1010011: c <= 9'b11100100;
				8'b1100001: c <= 9'b100100010;
				8'b110101: c <= 9'b110001000;
				8'b1000100: c <= 9'b11001011;
				8'b1010001: c <= 9'b110000010;
				8'b1010100: c <= 9'b10110110;
				8'b1100110: c <= 9'b101111010;
				8'b101010: c <= 9'b11001101;
				8'b1011110: c <= 9'b10111000;
				8'b1100111: c <= 9'b11110101;
				8'b1011010: c <= 9'b100110111;
				8'b1000010: c <= 9'b1111;
				8'b111101: c <= 9'b111000010;
				8'b110000: c <= 9'b10101110;
				8'b111110: c <= 9'b11111101;
				8'b1100010: c <= 9'b11110000;
				8'b1110000: c <= 9'b1110101;
				8'b1101001: c <= 9'b10101011;
				8'b1110011: c <= 9'b101001011;
				8'b1001100: c <= 9'b11101101;
				8'b100001: c <= 9'b10010000;
				8'b1000110: c <= 9'b1100;
				8'b1110010: c <= 9'b111011001;
				8'b1010000: c <= 9'b1100111;
				8'b1111010: c <= 9'b101100110;
				8'b1010101: c <= 9'b11111101;
				8'b111011: c <= 9'b101010011;
				8'b1001101: c <= 9'b10110001;
				8'b111111: c <= 9'b1010011;
				8'b1101110: c <= 9'b100100001;
				8'b1111011: c <= 9'b11111;
				8'b1001011: c <= 9'b1100;
				8'b1101111: c <= 9'b11000;
				8'b1101000: c <= 9'b1110111;
				8'b101100: c <= 9'b11011011;
				8'b100100: c <= 9'b110010101;
				8'b1111000: c <= 9'b111010000;
				8'b1000101: c <= 9'b1011110;
				8'b1011001: c <= 9'b100111101;
				8'b110100: c <= 9'b100001;
				8'b1111001: c <= 9'b101110111;
				8'b1110001: c <= 9'b100110;
				8'b1001111: c <= 9'b110101110;
				8'b1100101: c <= 9'b101010001;
				8'b1111110: c <= 9'b100010111;
				8'b1111100: c <= 9'b11011110;
				8'b1010110: c <= 9'b10001001;
				8'b110010: c <= 9'b101100101;
				8'b1101101: c <= 9'b101010100;
				8'b100011: c <= 9'b110110000;
				8'b1110101: c <= 9'b1100001;
				8'b1111101: c <= 9'b100111110;
				8'b101001: c <= 9'b110000000;
				8'b1010010: c <= 9'b1001111;
				8'b1011000: c <= 9'b10001011;
				8'b101110: c <= 9'b110001100;
				8'b1000001: c <= 9'b11111101;
				default: c <= 9'b0;
			endcase
			9'b10101110 : case(di)
				8'b1000011: c <= 9'b100010010;
				8'b101000: c <= 9'b10111;
				8'b111010: c <= 9'b11111000;
				8'b110110: c <= 9'b11010;
				8'b1100100: c <= 9'b100000000;
				8'b1000000: c <= 9'b100000100;
				8'b1110110: c <= 9'b111101111;
				8'b100101: c <= 9'b101010011;
				8'b101111: c <= 9'b110000101;
				8'b100110: c <= 9'b100011001;
				8'b1100011: c <= 9'b100010000;
				8'b1001000: c <= 9'b111110000;
				8'b111000: c <= 9'b110010100;
				8'b110001: c <= 9'b10;
				8'b1010111: c <= 9'b101010100;
				8'b1001110: c <= 9'b11001100;
				8'b1101010: c <= 9'b11100101;
				8'b1001001: c <= 9'b111100001;
				8'b1100000: c <= 9'b11000;
				8'b110111: c <= 9'b10101010;
				8'b1011101: c <= 9'b1111010;
				8'b1011011: c <= 9'b101101111;
				8'b111001: c <= 9'b110110110;
				8'b1001010: c <= 9'b101011111;
				8'b110011: c <= 9'b10011101;
				8'b1101100: c <= 9'b101100001;
				8'b1110111: c <= 9'b110000001;
				8'b101011: c <= 9'b101001010;
				8'b1101011: c <= 9'b10011010;
				8'b111100: c <= 9'b1000;
				8'b1000111: c <= 9'b101110010;
				8'b1011111: c <= 9'b1010110;
				8'b1110100: c <= 9'b10100011;
				8'b101101: c <= 9'b11110011;
				8'b1010011: c <= 9'b11010011;
				8'b1100001: c <= 9'b110000111;
				8'b110101: c <= 9'b101111001;
				8'b1000100: c <= 9'b10011100;
				8'b1010001: c <= 9'b10010101;
				8'b1010100: c <= 9'b1011100;
				8'b1100110: c <= 9'b101101011;
				8'b101010: c <= 9'b11010100;
				8'b1011110: c <= 9'b11001010;
				8'b1100111: c <= 9'b10101110;
				8'b1011010: c <= 9'b101110;
				8'b1000010: c <= 9'b10010011;
				8'b111101: c <= 9'b111100110;
				8'b110000: c <= 9'b101001000;
				8'b111110: c <= 9'b101110;
				8'b1100010: c <= 9'b100011101;
				8'b1110000: c <= 9'b111101001;
				8'b1101001: c <= 9'b1011001;
				8'b1110011: c <= 9'b100010010;
				8'b1001100: c <= 9'b10010000;
				8'b100001: c <= 9'b11101011;
				8'b1000110: c <= 9'b11110110;
				8'b1110010: c <= 9'b101100110;
				8'b1010000: c <= 9'b101101000;
				8'b1111010: c <= 9'b1010110;
				8'b1010101: c <= 9'b110000;
				8'b111011: c <= 9'b10111111;
				8'b1001101: c <= 9'b1011001;
				8'b111111: c <= 9'b11101001;
				8'b1101110: c <= 9'b10101100;
				8'b1111011: c <= 9'b110101001;
				8'b1001011: c <= 9'b11110101;
				8'b1101111: c <= 9'b101101100;
				8'b1101000: c <= 9'b11101000;
				8'b101100: c <= 9'b111111101;
				8'b100100: c <= 9'b11101;
				8'b1111000: c <= 9'b100000010;
				8'b1000101: c <= 9'b10100;
				8'b1011001: c <= 9'b10101100;
				8'b110100: c <= 9'b111011001;
				8'b1111001: c <= 9'b1101110;
				8'b1110001: c <= 9'b11111110;
				8'b1001111: c <= 9'b11111000;
				8'b1100101: c <= 9'b11011010;
				8'b1111110: c <= 9'b10101110;
				8'b1111100: c <= 9'b101100101;
				8'b1010110: c <= 9'b101110001;
				8'b110010: c <= 9'b101001001;
				8'b1101101: c <= 9'b110010;
				8'b100011: c <= 9'b10110110;
				8'b1110101: c <= 9'b10010011;
				8'b1111101: c <= 9'b1110000;
				8'b101001: c <= 9'b1100000;
				8'b1010010: c <= 9'b110011011;
				8'b1011000: c <= 9'b101010011;
				8'b101110: c <= 9'b10001100;
				8'b1000001: c <= 9'b100111011;
				default: c <= 9'b0;
			endcase
			9'b1000110 : case(di)
				8'b1000011: c <= 9'b1111011;
				8'b101000: c <= 9'b1000101;
				8'b111010: c <= 9'b1001111;
				8'b110110: c <= 9'b111001010;
				8'b1100100: c <= 9'b101000010;
				8'b1000000: c <= 9'b11110000;
				8'b1110110: c <= 9'b111000010;
				8'b100101: c <= 9'b10011000;
				8'b101111: c <= 9'b1;
				8'b100110: c <= 9'b101111010;
				8'b1100011: c <= 9'b10000101;
				8'b1001000: c <= 9'b110110;
				8'b111000: c <= 9'b100011000;
				8'b110001: c <= 9'b100011011;
				8'b1010111: c <= 9'b1100010;
				8'b1001110: c <= 9'b101111010;
				8'b1101010: c <= 9'b100011111;
				8'b1001001: c <= 9'b110100000;
				8'b1100000: c <= 9'b111111011;
				8'b110111: c <= 9'b100100000;
				8'b1011101: c <= 9'b10000111;
				8'b1011011: c <= 9'b10000101;
				8'b111001: c <= 9'b11011011;
				8'b1001010: c <= 9'b11100010;
				8'b110011: c <= 9'b10010;
				8'b1101100: c <= 9'b100100011;
				8'b1110111: c <= 9'b101100011;
				8'b101011: c <= 9'b101100100;
				8'b1101011: c <= 9'b100000001;
				8'b111100: c <= 9'b11111000;
				8'b1000111: c <= 9'b10001000;
				8'b1011111: c <= 9'b110100110;
				8'b1110100: c <= 9'b100110;
				8'b101101: c <= 9'b11001100;
				8'b1010011: c <= 9'b1011111;
				8'b1100001: c <= 9'b100010010;
				8'b110101: c <= 9'b110111010;
				8'b1000100: c <= 9'b100100001;
				8'b1010001: c <= 9'b110010101;
				8'b1010100: c <= 9'b101011011;
				8'b1100110: c <= 9'b100100101;
				8'b101010: c <= 9'b11010001;
				8'b1011110: c <= 9'b1010110;
				8'b1100111: c <= 9'b1101000;
				8'b1011010: c <= 9'b101100101;
				8'b1000010: c <= 9'b110110000;
				8'b111101: c <= 9'b101011110;
				8'b110000: c <= 9'b10100100;
				8'b111110: c <= 9'b10001110;
				8'b1100010: c <= 9'b1100010;
				8'b1110000: c <= 9'b110110011;
				8'b1101001: c <= 9'b110110100;
				8'b1110011: c <= 9'b11101111;
				8'b1001100: c <= 9'b100010110;
				8'b100001: c <= 9'b11100;
				8'b1000110: c <= 9'b101101000;
				8'b1110010: c <= 9'b100010100;
				8'b1010000: c <= 9'b10100000;
				8'b1111010: c <= 9'b100100111;
				8'b1010101: c <= 9'b110111110;
				8'b111011: c <= 9'b1111111;
				8'b1001101: c <= 9'b100011101;
				8'b111111: c <= 9'b101110100;
				8'b1101110: c <= 9'b111011011;
				8'b1111011: c <= 9'b110000110;
				8'b1001011: c <= 9'b100100110;
				8'b1101111: c <= 9'b10011;
				8'b1101000: c <= 9'b1100101;
				8'b101100: c <= 9'b11101000;
				8'b100100: c <= 9'b101100110;
				8'b1111000: c <= 9'b11010101;
				8'b1000101: c <= 9'b101100001;
				8'b1011001: c <= 9'b100010110;
				8'b110100: c <= 9'b100010101;
				8'b1111001: c <= 9'b1000011;
				8'b1110001: c <= 9'b101111010;
				8'b1001111: c <= 9'b1111000;
				8'b1100101: c <= 9'b10110100;
				8'b1111110: c <= 9'b10110011;
				8'b1111100: c <= 9'b110101110;
				8'b1010110: c <= 9'b100011100;
				8'b110010: c <= 9'b110001010;
				8'b1101101: c <= 9'b111111000;
				8'b100011: c <= 9'b111010111;
				8'b1110101: c <= 9'b1000011;
				8'b1111101: c <= 9'b1010011;
				8'b101001: c <= 9'b111100111;
				8'b1010010: c <= 9'b111101;
				8'b1011000: c <= 9'b11101100;
				8'b101110: c <= 9'b110010110;
				8'b1000001: c <= 9'b1000110;
				default: c <= 9'b0;
			endcase
			9'b1100101 : case(di)
				8'b1000011: c <= 9'b100010001;
				8'b101000: c <= 9'b10110;
				8'b111010: c <= 9'b10000;
				8'b110110: c <= 9'b111110011;
				8'b1100100: c <= 9'b100111011;
				8'b1000000: c <= 9'b100111010;
				8'b1110110: c <= 9'b1101111;
				8'b100101: c <= 9'b100101111;
				8'b101111: c <= 9'b100111000;
				8'b100110: c <= 9'b11;
				8'b1100011: c <= 9'b110110000;
				8'b1001000: c <= 9'b11110000;
				8'b111000: c <= 9'b101000101;
				8'b110001: c <= 9'b1110001;
				8'b1010111: c <= 9'b110011111;
				8'b1001110: c <= 9'b100111011;
				8'b1101010: c <= 9'b1101000;
				8'b1001001: c <= 9'b11100101;
				8'b1100000: c <= 9'b101010100;
				8'b110111: c <= 9'b1001;
				8'b1011101: c <= 9'b10011111;
				8'b1011011: c <= 9'b111001;
				8'b111001: c <= 9'b1000110;
				8'b1001010: c <= 9'b100111111;
				8'b110011: c <= 9'b100000110;
				8'b1101100: c <= 9'b111000;
				8'b1110111: c <= 9'b11101101;
				8'b101011: c <= 9'b100000000;
				8'b1101011: c <= 9'b100000100;
				8'b111100: c <= 9'b100110000;
				8'b1000111: c <= 9'b100001011;
				8'b1011111: c <= 9'b101011011;
				8'b1110100: c <= 9'b111001101;
				8'b101101: c <= 9'b111010000;
				8'b1010011: c <= 9'b10010000;
				8'b1100001: c <= 9'b1011010;
				8'b110101: c <= 9'b1011001;
				8'b1000100: c <= 9'b110010100;
				8'b1010001: c <= 9'b110011001;
				8'b1010100: c <= 9'b100011001;
				8'b1100110: c <= 9'b100100;
				8'b101010: c <= 9'b110011000;
				8'b1011110: c <= 9'b111001111;
				8'b1100111: c <= 9'b1010011;
				8'b1011010: c <= 9'b10110001;
				8'b1000010: c <= 9'b111100010;
				8'b111101: c <= 9'b101101010;
				8'b110000: c <= 9'b11110101;
				8'b111110: c <= 9'b11010100;
				8'b1100010: c <= 9'b101001010;
				8'b1110000: c <= 9'b1011001;
				8'b1101001: c <= 9'b10000000;
				8'b1110011: c <= 9'b101100110;
				8'b1001100: c <= 9'b100000001;
				8'b100001: c <= 9'b101001000;
				8'b1000110: c <= 9'b10001100;
				8'b1110010: c <= 9'b10111101;
				8'b1010000: c <= 9'b101011011;
				8'b1111010: c <= 9'b100101000;
				8'b1010101: c <= 9'b111100001;
				8'b111011: c <= 9'b100011100;
				8'b1001101: c <= 9'b100111110;
				8'b111111: c <= 9'b111100010;
				8'b1101110: c <= 9'b111101010;
				8'b1111011: c <= 9'b111101;
				8'b1001011: c <= 9'b10010110;
				8'b1101111: c <= 9'b10001101;
				8'b1101000: c <= 9'b111110011;
				8'b101100: c <= 9'b1100100;
				8'b100100: c <= 9'b100001111;
				8'b1111000: c <= 9'b110001111;
				8'b1000101: c <= 9'b10111110;
				8'b1011001: c <= 9'b101101001;
				8'b110100: c <= 9'b11011;
				8'b1111001: c <= 9'b101110100;
				8'b1110001: c <= 9'b1111110;
				8'b1001111: c <= 9'b10;
				8'b1100101: c <= 9'b110100110;
				8'b1111110: c <= 9'b111011101;
				8'b1111100: c <= 9'b1011001;
				8'b1010110: c <= 9'b1000101;
				8'b110010: c <= 9'b100001111;
				8'b1101101: c <= 9'b110100;
				8'b100011: c <= 9'b101111000;
				8'b1110101: c <= 9'b10111010;
				8'b1111101: c <= 9'b11000011;
				8'b101001: c <= 9'b110011100;
				8'b1010010: c <= 9'b110101111;
				8'b1011000: c <= 9'b11001001;
				8'b101110: c <= 9'b101111111;
				8'b1000001: c <= 9'b1011000;
				default: c <= 9'b0;
			endcase
			9'b101011000 : case(di)
				8'b1000011: c <= 9'b111010100;
				8'b101000: c <= 9'b11000;
				8'b111010: c <= 9'b100100001;
				8'b110110: c <= 9'b100011100;
				8'b1100100: c <= 9'b11011;
				8'b1000000: c <= 9'b101010001;
				8'b1110110: c <= 9'b111110110;
				8'b100101: c <= 9'b100110010;
				8'b101111: c <= 9'b1010011;
				8'b100110: c <= 9'b101101011;
				8'b1100011: c <= 9'b101001111;
				8'b1001000: c <= 9'b11101;
				8'b111000: c <= 9'b100110011;
				8'b110001: c <= 9'b11011110;
				8'b1010111: c <= 9'b1011;
				8'b1001110: c <= 9'b100101001;
				8'b1101010: c <= 9'b111101000;
				8'b1001001: c <= 9'b101000010;
				8'b1100000: c <= 9'b111100010;
				8'b110111: c <= 9'b1010011;
				8'b1011101: c <= 9'b101011101;
				8'b1011011: c <= 9'b1101000;
				8'b111001: c <= 9'b111110001;
				8'b1001010: c <= 9'b100101000;
				8'b110011: c <= 9'b100100;
				8'b1101100: c <= 9'b1000101;
				8'b1110111: c <= 9'b1011110;
				8'b101011: c <= 9'b10001000;
				8'b1101011: c <= 9'b1010011;
				8'b111100: c <= 9'b1000000;
				8'b1000111: c <= 9'b111001111;
				8'b1011111: c <= 9'b1001110;
				8'b1110100: c <= 9'b10110010;
				8'b101101: c <= 9'b110000010;
				8'b1010011: c <= 9'b1100100;
				8'b1100001: c <= 9'b110011011;
				8'b110101: c <= 9'b10101011;
				8'b1000100: c <= 9'b111100101;
				8'b1010001: c <= 9'b11100010;
				8'b1010100: c <= 9'b111100;
				8'b1100110: c <= 9'b101011;
				8'b101010: c <= 9'b100000101;
				8'b1011110: c <= 9'b100101001;
				8'b1100111: c <= 9'b101111110;
				8'b1011010: c <= 9'b101001010;
				8'b1000010: c <= 9'b1101101;
				8'b111101: c <= 9'b101001110;
				8'b110000: c <= 9'b111001010;
				8'b111110: c <= 9'b111100111;
				8'b1100010: c <= 9'b11111010;
				8'b1110000: c <= 9'b1000000;
				8'b1101001: c <= 9'b1100;
				8'b1110011: c <= 9'b111100110;
				8'b1001100: c <= 9'b1;
				8'b100001: c <= 9'b101001010;
				8'b1000110: c <= 9'b10110001;
				8'b1110010: c <= 9'b111101110;
				8'b1010000: c <= 9'b101100011;
				8'b1111010: c <= 9'b111001;
				8'b1010101: c <= 9'b11001110;
				8'b111011: c <= 9'b10111100;
				8'b1001101: c <= 9'b110001100;
				8'b111111: c <= 9'b100100;
				8'b1101110: c <= 9'b101001011;
				8'b1111011: c <= 9'b111110110;
				8'b1001011: c <= 9'b100001;
				8'b1101111: c <= 9'b11111010;
				8'b1101000: c <= 9'b100101001;
				8'b101100: c <= 9'b11100111;
				8'b100100: c <= 9'b101100;
				8'b1111000: c <= 9'b10100011;
				8'b1000101: c <= 9'b111100100;
				8'b1011001: c <= 9'b110011111;
				8'b110100: c <= 9'b11001001;
				8'b1111001: c <= 9'b101000101;
				8'b1110001: c <= 9'b11010001;
				8'b1001111: c <= 9'b111111111;
				8'b1100101: c <= 9'b111010110;
				8'b1111110: c <= 9'b1101110;
				8'b1111100: c <= 9'b110100110;
				8'b1010110: c <= 9'b11001101;
				8'b110010: c <= 9'b100100;
				8'b1101101: c <= 9'b111111;
				8'b100011: c <= 9'b100011001;
				8'b1110101: c <= 9'b1001111;
				8'b1111101: c <= 9'b1000010;
				8'b101001: c <= 9'b10001110;
				8'b1010010: c <= 9'b100000001;
				8'b1011000: c <= 9'b10001001;
				8'b101110: c <= 9'b110110111;
				8'b1000001: c <= 9'b101011111;
				default: c <= 9'b0;
			endcase
			9'b110110100 : case(di)
				8'b1000011: c <= 9'b11110001;
				8'b101000: c <= 9'b111111111;
				8'b111010: c <= 9'b11001000;
				8'b110110: c <= 9'b11111001;
				8'b1100100: c <= 9'b11100111;
				8'b1000000: c <= 9'b11100001;
				8'b1110110: c <= 9'b101110010;
				8'b100101: c <= 9'b10000;
				8'b101111: c <= 9'b10011000;
				8'b100110: c <= 9'b1000001;
				8'b1100011: c <= 9'b111101110;
				8'b1001000: c <= 9'b101000011;
				8'b111000: c <= 9'b110001011;
				8'b110001: c <= 9'b101011101;
				8'b1010111: c <= 9'b1110001;
				8'b1001110: c <= 9'b1100010;
				8'b1101010: c <= 9'b1101010;
				8'b1001001: c <= 9'b100011;
				8'b1100000: c <= 9'b100011010;
				8'b110111: c <= 9'b101110010;
				8'b1011101: c <= 9'b11010101;
				8'b1011011: c <= 9'b1100010;
				8'b111001: c <= 9'b110011000;
				8'b1001010: c <= 9'b110010100;
				8'b110011: c <= 9'b1100111;
				8'b1101100: c <= 9'b101100100;
				8'b1110111: c <= 9'b11011110;
				8'b101011: c <= 9'b10001110;
				8'b1101011: c <= 9'b110101111;
				8'b111100: c <= 9'b11100001;
				8'b1000111: c <= 9'b11000100;
				8'b1011111: c <= 9'b110110;
				8'b1110100: c <= 9'b1011000;
				8'b101101: c <= 9'b101001001;
				8'b1010011: c <= 9'b111110101;
				8'b1100001: c <= 9'b1010001;
				8'b110101: c <= 9'b101110100;
				8'b1000100: c <= 9'b1011;
				8'b1010001: c <= 9'b1011;
				8'b1010100: c <= 9'b100011001;
				8'b1100110: c <= 9'b111101;
				8'b101010: c <= 9'b111011111;
				8'b1011110: c <= 9'b101011010;
				8'b1100111: c <= 9'b111010001;
				8'b1011010: c <= 9'b111101110;
				8'b1000010: c <= 9'b110110000;
				8'b111101: c <= 9'b100001100;
				8'b110000: c <= 9'b1110101;
				8'b111110: c <= 9'b110000010;
				8'b1100010: c <= 9'b11010001;
				8'b1110000: c <= 9'b101000001;
				8'b1101001: c <= 9'b110111011;
				8'b1110011: c <= 9'b111101;
				8'b1001100: c <= 9'b10010000;
				8'b100001: c <= 9'b101111110;
				8'b1000110: c <= 9'b1100010;
				8'b1110010: c <= 9'b101100001;
				8'b1010000: c <= 9'b110101111;
				8'b1111010: c <= 9'b100100;
				8'b1010101: c <= 9'b1111001;
				8'b111011: c <= 9'b111011;
				8'b1001101: c <= 9'b11111110;
				8'b111111: c <= 9'b11101;
				8'b1101110: c <= 9'b100000101;
				8'b1111011: c <= 9'b101011;
				8'b1001011: c <= 9'b11001000;
				8'b1101111: c <= 9'b11111110;
				8'b1101000: c <= 9'b10101000;
				8'b101100: c <= 9'b11101101;
				8'b100100: c <= 9'b111111011;
				8'b1111000: c <= 9'b111;
				8'b1000101: c <= 9'b11100010;
				8'b1011001: c <= 9'b11111001;
				8'b110100: c <= 9'b100011010;
				8'b1111001: c <= 9'b11110011;
				8'b1110001: c <= 9'b111;
				8'b1001111: c <= 9'b110001101;
				8'b1100101: c <= 9'b11001001;
				8'b1111110: c <= 9'b111100110;
				8'b1111100: c <= 9'b110;
				8'b1010110: c <= 9'b111100011;
				8'b110010: c <= 9'b110101101;
				8'b1101101: c <= 9'b100110100;
				8'b100011: c <= 9'b10001001;
				8'b1110101: c <= 9'b100110110;
				8'b1111101: c <= 9'b100100001;
				8'b101001: c <= 9'b10001110;
				8'b1010010: c <= 9'b110001011;
				8'b1011000: c <= 9'b11011;
				8'b101110: c <= 9'b111001110;
				8'b1000001: c <= 9'b11111001;
				default: c <= 9'b0;
			endcase
			9'b11010001 : case(di)
				8'b1000011: c <= 9'b101010100;
				8'b101000: c <= 9'b101111001;
				8'b111010: c <= 9'b11111110;
				8'b110110: c <= 9'b101101110;
				8'b1100100: c <= 9'b10110010;
				8'b1000000: c <= 9'b1011;
				8'b1110110: c <= 9'b100100111;
				8'b100101: c <= 9'b110001;
				8'b101111: c <= 9'b101000111;
				8'b100110: c <= 9'b11000111;
				8'b1100011: c <= 9'b11101111;
				8'b1001000: c <= 9'b111100;
				8'b111000: c <= 9'b1;
				8'b110001: c <= 9'b101110;
				8'b1010111: c <= 9'b11100111;
				8'b1001110: c <= 9'b110100110;
				8'b1101010: c <= 9'b110111110;
				8'b1001001: c <= 9'b1011011;
				8'b1100000: c <= 9'b11100110;
				8'b110111: c <= 9'b1101101;
				8'b1011101: c <= 9'b11100110;
				8'b1011011: c <= 9'b101001001;
				8'b111001: c <= 9'b10001000;
				8'b1001010: c <= 9'b100001001;
				8'b110011: c <= 9'b10010001;
				8'b1101100: c <= 9'b110011100;
				8'b1110111: c <= 9'b10101000;
				8'b101011: c <= 9'b11110000;
				8'b1101011: c <= 9'b100111001;
				8'b111100: c <= 9'b11100011;
				8'b1000111: c <= 9'b111001110;
				8'b1011111: c <= 9'b110010001;
				8'b1110100: c <= 9'b101101011;
				8'b101101: c <= 9'b111010001;
				8'b1010011: c <= 9'b100010011;
				8'b1100001: c <= 9'b100101101;
				8'b110101: c <= 9'b100101;
				8'b1000100: c <= 9'b101100010;
				8'b1010001: c <= 9'b10000101;
				8'b1010100: c <= 9'b110011000;
				8'b1100110: c <= 9'b101100001;
				8'b101010: c <= 9'b110111010;
				8'b1011110: c <= 9'b111111111;
				8'b1100111: c <= 9'b1010011;
				8'b1011010: c <= 9'b10000000;
				8'b1000010: c <= 9'b100001101;
				8'b111101: c <= 9'b111101100;
				8'b110000: c <= 9'b101010000;
				8'b111110: c <= 9'b110111010;
				8'b1100010: c <= 9'b100100011;
				8'b1110000: c <= 9'b101100011;
				8'b1101001: c <= 9'b100001;
				8'b1110011: c <= 9'b110111100;
				8'b1001100: c <= 9'b11000011;
				8'b100001: c <= 9'b11010010;
				8'b1000110: c <= 9'b111111111;
				8'b1110010: c <= 9'b100011001;
				8'b1010000: c <= 9'b1000110;
				8'b1111010: c <= 9'b1101101;
				8'b1010101: c <= 9'b11010001;
				8'b111011: c <= 9'b11010;
				8'b1001101: c <= 9'b1011110;
				8'b111111: c <= 9'b1100010;
				8'b1101110: c <= 9'b10111001;
				8'b1111011: c <= 9'b110010011;
				8'b1001011: c <= 9'b110000110;
				8'b1101111: c <= 9'b110111010;
				8'b1101000: c <= 9'b111110101;
				8'b101100: c <= 9'b101010001;
				8'b100100: c <= 9'b110001111;
				8'b1111000: c <= 9'b100111010;
				8'b1000101: c <= 9'b1111101;
				8'b1011001: c <= 9'b1011100;
				8'b110100: c <= 9'b11111110;
				8'b1111001: c <= 9'b100001110;
				8'b1110001: c <= 9'b1111110;
				8'b1001111: c <= 9'b10100100;
				8'b1100101: c <= 9'b111011010;
				8'b1111110: c <= 9'b110100000;
				8'b1111100: c <= 9'b100000111;
				8'b1010110: c <= 9'b110011011;
				8'b110010: c <= 9'b101101010;
				8'b1101101: c <= 9'b1000011;
				8'b100011: c <= 9'b10101010;
				8'b1110101: c <= 9'b110011;
				8'b1111101: c <= 9'b111010000;
				8'b101001: c <= 9'b11000111;
				8'b1010010: c <= 9'b111100100;
				8'b1011000: c <= 9'b101000101;
				8'b101110: c <= 9'b10110;
				8'b1000001: c <= 9'b110000010;
				default: c <= 9'b0;
			endcase
			9'b111100100 : case(di)
				8'b1000011: c <= 9'b100010;
				8'b101000: c <= 9'b101011011;
				8'b111010: c <= 9'b10000101;
				8'b110110: c <= 9'b110111111;
				8'b1100100: c <= 9'b100000101;
				8'b1000000: c <= 9'b11111;
				8'b1110110: c <= 9'b111010110;
				8'b100101: c <= 9'b10001011;
				8'b101111: c <= 9'b110010010;
				8'b100110: c <= 9'b110010001;
				8'b1100011: c <= 9'b111100110;
				8'b1001000: c <= 9'b1111101;
				8'b111000: c <= 9'b101101001;
				8'b110001: c <= 9'b111000011;
				8'b1010111: c <= 9'b100111;
				8'b1001110: c <= 9'b1011;
				8'b1101010: c <= 9'b101010101;
				8'b1001001: c <= 9'b10011111;
				8'b1100000: c <= 9'b11000;
				8'b110111: c <= 9'b1100111;
				8'b1011101: c <= 9'b11010000;
				8'b1011011: c <= 9'b11011010;
				8'b111001: c <= 9'b101110101;
				8'b1001010: c <= 9'b111010111;
				8'b110011: c <= 9'b110110111;
				8'b1101100: c <= 9'b100010111;
				8'b1110111: c <= 9'b11001111;
				8'b101011: c <= 9'b101000010;
				8'b1101011: c <= 9'b101101100;
				8'b111100: c <= 9'b11;
				8'b1000111: c <= 9'b100;
				8'b1011111: c <= 9'b11111011;
				8'b1110100: c <= 9'b10101000;
				8'b101101: c <= 9'b111111011;
				8'b1010011: c <= 9'b1110;
				8'b1100001: c <= 9'b10100011;
				8'b110101: c <= 9'b101001;
				8'b1000100: c <= 9'b10010101;
				8'b1010001: c <= 9'b110100111;
				8'b1010100: c <= 9'b11;
				8'b1100110: c <= 9'b101110011;
				8'b101010: c <= 9'b10;
				8'b1011110: c <= 9'b11111000;
				8'b1100111: c <= 9'b100010111;
				8'b1011010: c <= 9'b11011011;
				8'b1000010: c <= 9'b1100;
				8'b111101: c <= 9'b11000110;
				8'b110000: c <= 9'b111010001;
				8'b111110: c <= 9'b11010111;
				8'b1100010: c <= 9'b11010000;
				8'b1110000: c <= 9'b1111000;
				8'b1101001: c <= 9'b11111011;
				8'b1110011: c <= 9'b101111001;
				8'b1001100: c <= 9'b10110110;
				8'b100001: c <= 9'b1011010;
				8'b1000110: c <= 9'b100000011;
				8'b1110010: c <= 9'b100110000;
				8'b1010000: c <= 9'b10000;
				8'b1111010: c <= 9'b111110101;
				8'b1010101: c <= 9'b11100111;
				8'b111011: c <= 9'b110011010;
				8'b1001101: c <= 9'b111110000;
				8'b111111: c <= 9'b111001;
				8'b1101110: c <= 9'b110001111;
				8'b1111011: c <= 9'b1010110;
				8'b1001011: c <= 9'b10101100;
				8'b1101111: c <= 9'b111111;
				8'b1101000: c <= 9'b10111011;
				8'b101100: c <= 9'b111010010;
				8'b100100: c <= 9'b100100111;
				8'b1111000: c <= 9'b110011100;
				8'b1000101: c <= 9'b100101110;
				8'b1011001: c <= 9'b1111;
				8'b110100: c <= 9'b10011010;
				8'b1111001: c <= 9'b1110;
				8'b1110001: c <= 9'b1001110;
				8'b1001111: c <= 9'b110111000;
				8'b1100101: c <= 9'b11110011;
				8'b1111110: c <= 9'b110000101;
				8'b1111100: c <= 9'b111000000;
				8'b1010110: c <= 9'b100111010;
				8'b110010: c <= 9'b110001111;
				8'b1101101: c <= 9'b100100101;
				8'b100011: c <= 9'b11010;
				8'b1110101: c <= 9'b1110011;
				8'b1111101: c <= 9'b101110010;
				8'b101001: c <= 9'b11011000;
				8'b1010010: c <= 9'b101101111;
				8'b1011000: c <= 9'b110111;
				8'b101110: c <= 9'b11101101;
				8'b1000001: c <= 9'b111001;
				default: c <= 9'b0;
			endcase
			9'b111110000 : case(di)
				8'b1000011: c <= 9'b111011100;
				8'b101000: c <= 9'b110100000;
				8'b111010: c <= 9'b111010001;
				8'b110110: c <= 9'b111001111;
				8'b1100100: c <= 9'b11001101;
				8'b1000000: c <= 9'b110;
				8'b1110110: c <= 9'b110010001;
				8'b100101: c <= 9'b11100;
				8'b101111: c <= 9'b1111000;
				8'b100110: c <= 9'b111111010;
				8'b1100011: c <= 9'b101011010;
				8'b1001000: c <= 9'b110011011;
				8'b111000: c <= 9'b1100110;
				8'b110001: c <= 9'b110011;
				8'b1010111: c <= 9'b110101;
				8'b1001110: c <= 9'b110000001;
				8'b1101010: c <= 9'b10101;
				8'b1001001: c <= 9'b111010100;
				8'b1100000: c <= 9'b1011001;
				8'b110111: c <= 9'b1111110;
				8'b1011101: c <= 9'b101010110;
				8'b1011011: c <= 9'b101101100;
				8'b111001: c <= 9'b101001110;
				8'b1001010: c <= 9'b101010100;
				8'b110011: c <= 9'b10000111;
				8'b1101100: c <= 9'b100100110;
				8'b1110111: c <= 9'b11110011;
				8'b101011: c <= 9'b11101;
				8'b1101011: c <= 9'b10101110;
				8'b111100: c <= 9'b111110110;
				8'b1000111: c <= 9'b100000101;
				8'b1011111: c <= 9'b100110;
				8'b1110100: c <= 9'b1011010;
				8'b101101: c <= 9'b10111;
				8'b1010011: c <= 9'b1000111;
				8'b1100001: c <= 9'b10110001;
				8'b110101: c <= 9'b100000001;
				8'b1000100: c <= 9'b10101101;
				8'b1010001: c <= 9'b11101100;
				8'b1010100: c <= 9'b10110110;
				8'b1100110: c <= 9'b101100;
				8'b101010: c <= 9'b1100000;
				8'b1011110: c <= 9'b101000111;
				8'b1100111: c <= 9'b11101111;
				8'b1011010: c <= 9'b111101001;
				8'b1000010: c <= 9'b110011001;
				8'b111101: c <= 9'b100011001;
				8'b110000: c <= 9'b10000101;
				8'b111110: c <= 9'b111001111;
				8'b1100010: c <= 9'b110010;
				8'b1110000: c <= 9'b10101001;
				8'b1101001: c <= 9'b1011000;
				8'b1110011: c <= 9'b111011101;
				8'b1001100: c <= 9'b11001110;
				8'b100001: c <= 9'b110001011;
				8'b1000110: c <= 9'b1101100;
				8'b1110010: c <= 9'b110011001;
				8'b1010000: c <= 9'b101000111;
				8'b1111010: c <= 9'b11001011;
				8'b1010101: c <= 9'b11001111;
				8'b111011: c <= 9'b110000101;
				8'b1001101: c <= 9'b100100;
				8'b111111: c <= 9'b110011000;
				8'b1101110: c <= 9'b100101100;
				8'b1111011: c <= 9'b110001001;
				8'b1001011: c <= 9'b1101100;
				8'b1101111: c <= 9'b111001011;
				8'b1101000: c <= 9'b10110101;
				8'b101100: c <= 9'b1101110;
				8'b100100: c <= 9'b10110011;
				8'b1111000: c <= 9'b1000111;
				8'b1000101: c <= 9'b10111;
				8'b1011001: c <= 9'b101111001;
				8'b110100: c <= 9'b10001101;
				8'b1111001: c <= 9'b101001;
				8'b1110001: c <= 9'b101000010;
				8'b1001111: c <= 9'b100111101;
				8'b1100101: c <= 9'b110111001;
				8'b1111110: c <= 9'b110100100;
				8'b1111100: c <= 9'b11101101;
				8'b1010110: c <= 9'b1111100;
				8'b110010: c <= 9'b110010111;
				8'b1101101: c <= 9'b110010111;
				8'b100011: c <= 9'b101001010;
				8'b1110101: c <= 9'b110001001;
				8'b1111101: c <= 9'b100000000;
				8'b101001: c <= 9'b110010111;
				8'b1010010: c <= 9'b10110100;
				8'b1011000: c <= 9'b10001010;
				8'b101110: c <= 9'b100000111;
				8'b1000001: c <= 9'b100000010;
				default: c <= 9'b0;
			endcase
			9'b1111011 : case(di)
				8'b1000011: c <= 9'b111110110;
				8'b101000: c <= 9'b101100101;
				8'b111010: c <= 9'b1001101;
				8'b110110: c <= 9'b11001010;
				8'b1100100: c <= 9'b101010101;
				8'b1000000: c <= 9'b1001;
				8'b1110110: c <= 9'b10100011;
				8'b100101: c <= 9'b1011100;
				8'b101111: c <= 9'b1100;
				8'b100110: c <= 9'b11110001;
				8'b1100011: c <= 9'b10001010;
				8'b1001000: c <= 9'b100101001;
				8'b111000: c <= 9'b11001100;
				8'b110001: c <= 9'b100111001;
				8'b1010111: c <= 9'b111100011;
				8'b1001110: c <= 9'b10111101;
				8'b1101010: c <= 9'b1110010;
				8'b1001001: c <= 9'b101010001;
				8'b1100000: c <= 9'b1000010;
				8'b110111: c <= 9'b10010;
				8'b1011101: c <= 9'b1111111;
				8'b1011011: c <= 9'b10000010;
				8'b111001: c <= 9'b10100011;
				8'b1001010: c <= 9'b11011;
				8'b110011: c <= 9'b11001010;
				8'b1101100: c <= 9'b11101101;
				8'b1110111: c <= 9'b10001011;
				8'b101011: c <= 9'b11;
				8'b1101011: c <= 9'b100001001;
				8'b111100: c <= 9'b11111110;
				8'b1000111: c <= 9'b1001010;
				8'b1011111: c <= 9'b1101000;
				8'b1110100: c <= 9'b100101;
				8'b101101: c <= 9'b111111001;
				8'b1010011: c <= 9'b1010011;
				8'b1100001: c <= 9'b10110110;
				8'b110101: c <= 9'b11100001;
				8'b1000100: c <= 9'b10011011;
				8'b1010001: c <= 9'b10000110;
				8'b1010100: c <= 9'b101000011;
				8'b1100110: c <= 9'b101100110;
				8'b101010: c <= 9'b101110110;
				8'b1011110: c <= 9'b10100111;
				8'b1100111: c <= 9'b100101110;
				8'b1011010: c <= 9'b10101010;
				8'b1000010: c <= 9'b11110110;
				8'b111101: c <= 9'b10101101;
				8'b110000: c <= 9'b11000001;
				8'b111110: c <= 9'b100011001;
				8'b1100010: c <= 9'b1111;
				8'b1110000: c <= 9'b10110;
				8'b1101001: c <= 9'b101010111;
				8'b1110011: c <= 9'b100111111;
				8'b1001100: c <= 9'b110011001;
				8'b100001: c <= 9'b110101110;
				8'b1000110: c <= 9'b11011000;
				8'b1110010: c <= 9'b11;
				8'b1010000: c <= 9'b1000110;
				8'b1111010: c <= 9'b11011000;
				8'b1010101: c <= 9'b11011100;
				8'b111011: c <= 9'b10110011;
				8'b1001101: c <= 9'b111011011;
				8'b111111: c <= 9'b11111011;
				8'b1101110: c <= 9'b101011110;
				8'b1111011: c <= 9'b110011001;
				8'b1001011: c <= 9'b101011010;
				8'b1101111: c <= 9'b110001001;
				8'b1101000: c <= 9'b1001100;
				8'b101100: c <= 9'b10110010;
				8'b100100: c <= 9'b111011111;
				8'b1111000: c <= 9'b100011001;
				8'b1000101: c <= 9'b10001100;
				8'b1011001: c <= 9'b110110100;
				8'b110100: c <= 9'b110010001;
				8'b1111001: c <= 9'b1100100;
				8'b1110001: c <= 9'b110011101;
				8'b1001111: c <= 9'b101010001;
				8'b1100101: c <= 9'b11100111;
				8'b1111110: c <= 9'b11100010;
				8'b1111100: c <= 9'b100010010;
				8'b1010110: c <= 9'b111111110;
				8'b110010: c <= 9'b101000010;
				8'b1101101: c <= 9'b110010001;
				8'b100011: c <= 9'b111101010;
				8'b1110101: c <= 9'b111011111;
				8'b1111101: c <= 9'b10101;
				8'b101001: c <= 9'b11011010;
				8'b1010010: c <= 9'b1000110;
				8'b1011000: c <= 9'b100100111;
				8'b101110: c <= 9'b10101101;
				8'b1000001: c <= 9'b1110011;
				default: c <= 9'b0;
			endcase
			9'b11110110 : case(di)
				8'b1000011: c <= 9'b110011100;
				8'b101000: c <= 9'b10001100;
				8'b111010: c <= 9'b111001;
				8'b110110: c <= 9'b111010111;
				8'b1100100: c <= 9'b111100001;
				8'b1000000: c <= 9'b1111110;
				8'b1110110: c <= 9'b10101001;
				8'b100101: c <= 9'b1;
				8'b101111: c <= 9'b11100000;
				8'b100110: c <= 9'b111010;
				8'b1100011: c <= 9'b1000000;
				8'b1001000: c <= 9'b110011010;
				8'b111000: c <= 9'b110101011;
				8'b110001: c <= 9'b110001111;
				8'b1010111: c <= 9'b110000110;
				8'b1001110: c <= 9'b10000001;
				8'b1101010: c <= 9'b110011010;
				8'b1001001: c <= 9'b100010010;
				8'b1100000: c <= 9'b100001;
				8'b110111: c <= 9'b11101101;
				8'b1011101: c <= 9'b110110100;
				8'b1011011: c <= 9'b11100;
				8'b111001: c <= 9'b111000100;
				8'b1001010: c <= 9'b110011100;
				8'b110011: c <= 9'b101100110;
				8'b1101100: c <= 9'b11100011;
				8'b1110111: c <= 9'b11101011;
				8'b101011: c <= 9'b1010111;
				8'b1101011: c <= 9'b100100101;
				8'b111100: c <= 9'b1101111;
				8'b1000111: c <= 9'b11111110;
				8'b1011111: c <= 9'b11010000;
				8'b1110100: c <= 9'b101101011;
				8'b101101: c <= 9'b110010011;
				8'b1010011: c <= 9'b111011010;
				8'b1100001: c <= 9'b1010111;
				8'b110101: c <= 9'b10100000;
				8'b1000100: c <= 9'b11001;
				8'b1010001: c <= 9'b1100010;
				8'b1010100: c <= 9'b110111110;
				8'b1100110: c <= 9'b110;
				8'b101010: c <= 9'b10011111;
				8'b1011110: c <= 9'b1001111;
				8'b1100111: c <= 9'b1110101;
				8'b1011010: c <= 9'b11101101;
				8'b1000010: c <= 9'b110000001;
				8'b111101: c <= 9'b101100010;
				8'b110000: c <= 9'b11100;
				8'b111110: c <= 9'b101000010;
				8'b1100010: c <= 9'b10011100;
				8'b1110000: c <= 9'b10111110;
				8'b1101001: c <= 9'b1001010;
				8'b1110011: c <= 9'b110011000;
				8'b1001100: c <= 9'b10000101;
				8'b100001: c <= 9'b1111101;
				8'b1000110: c <= 9'b10111001;
				8'b1110010: c <= 9'b110101110;
				8'b1010000: c <= 9'b11000010;
				8'b1111010: c <= 9'b111100;
				8'b1010101: c <= 9'b111111;
				8'b111011: c <= 9'b110100000;
				8'b1001101: c <= 9'b1111010;
				8'b111111: c <= 9'b101110111;
				8'b1101110: c <= 9'b111110000;
				8'b1111011: c <= 9'b111011;
				8'b1001011: c <= 9'b110100011;
				8'b1101111: c <= 9'b111;
				8'b1101000: c <= 9'b101000110;
				8'b101100: c <= 9'b11110110;
				8'b100100: c <= 9'b111010110;
				8'b1111000: c <= 9'b10110001;
				8'b1000101: c <= 9'b10000;
				8'b1011001: c <= 9'b110100110;
				8'b110100: c <= 9'b1011000;
				8'b1111001: c <= 9'b1101;
				8'b1110001: c <= 9'b11111001;
				8'b1001111: c <= 9'b111000010;
				8'b1100101: c <= 9'b1101010;
				8'b1111110: c <= 9'b10000011;
				8'b1111100: c <= 9'b11001111;
				8'b1010110: c <= 9'b10011111;
				8'b110010: c <= 9'b100011010;
				8'b1101101: c <= 9'b101101111;
				8'b100011: c <= 9'b10111000;
				8'b1110101: c <= 9'b10010000;
				8'b1111101: c <= 9'b110010100;
				8'b101001: c <= 9'b1010111;
				8'b1010010: c <= 9'b100101111;
				8'b1011000: c <= 9'b100000110;
				8'b101110: c <= 9'b10111110;
				8'b1000001: c <= 9'b11000100;
				default: c <= 9'b0;
			endcase
			9'b100011 : case(di)
				8'b1000011: c <= 9'b11000011;
				8'b101000: c <= 9'b101011010;
				8'b111010: c <= 9'b110110100;
				8'b110110: c <= 9'b110110110;
				8'b1100100: c <= 9'b101101101;
				8'b1000000: c <= 9'b110001000;
				8'b1110110: c <= 9'b1100110;
				8'b100101: c <= 9'b11001010;
				8'b101111: c <= 9'b1010011;
				8'b100110: c <= 9'b111111101;
				8'b1100011: c <= 9'b11011010;
				8'b1001000: c <= 9'b10101010;
				8'b111000: c <= 9'b10111011;
				8'b110001: c <= 9'b101001111;
				8'b1010111: c <= 9'b100010001;
				8'b1001110: c <= 9'b1111100;
				8'b1101010: c <= 9'b110110010;
				8'b1001001: c <= 9'b1000101;
				8'b1100000: c <= 9'b11110000;
				8'b110111: c <= 9'b110000;
				8'b1011101: c <= 9'b100010011;
				8'b1011011: c <= 9'b101101100;
				8'b111001: c <= 9'b11000011;
				8'b1001010: c <= 9'b10010110;
				8'b110011: c <= 9'b1001101;
				8'b1101100: c <= 9'b110000;
				8'b1110111: c <= 9'b11111110;
				8'b101011: c <= 9'b11101011;
				8'b1101011: c <= 9'b10001110;
				8'b111100: c <= 9'b10100000;
				8'b1000111: c <= 9'b100100;
				8'b1011111: c <= 9'b11101001;
				8'b1110100: c <= 9'b1111010;
				8'b101101: c <= 9'b100011101;
				8'b1010011: c <= 9'b110000101;
				8'b1100001: c <= 9'b111011011;
				8'b110101: c <= 9'b110001001;
				8'b1000100: c <= 9'b10110110;
				8'b1010001: c <= 9'b10010001;
				8'b1010100: c <= 9'b10000110;
				8'b1100110: c <= 9'b1011000;
				8'b101010: c <= 9'b1110101;
				8'b1011110: c <= 9'b111100110;
				8'b1100111: c <= 9'b11001111;
				8'b1011010: c <= 9'b1010001;
				8'b1000010: c <= 9'b10011111;
				8'b111101: c <= 9'b111101111;
				8'b110000: c <= 9'b110000110;
				8'b111110: c <= 9'b11001;
				8'b1100010: c <= 9'b101101001;
				8'b1110000: c <= 9'b1000110;
				8'b1101001: c <= 9'b10110010;
				8'b1110011: c <= 9'b1010101;
				8'b1001100: c <= 9'b100101110;
				8'b100001: c <= 9'b1100000;
				8'b1000110: c <= 9'b1110111;
				8'b1110010: c <= 9'b100001010;
				8'b1010000: c <= 9'b1000000;
				8'b1111010: c <= 9'b100101011;
				8'b1010101: c <= 9'b110111010;
				8'b111011: c <= 9'b10000;
				8'b1001101: c <= 9'b1101101;
				8'b111111: c <= 9'b111111011;
				8'b1101110: c <= 9'b11111101;
				8'b1111011: c <= 9'b1110000;
				8'b1001011: c <= 9'b11011000;
				8'b1101111: c <= 9'b10000010;
				8'b1101000: c <= 9'b111011110;
				8'b101100: c <= 9'b1011100;
				8'b100100: c <= 9'b100101000;
				8'b1111000: c <= 9'b110011110;
				8'b1000101: c <= 9'b11101000;
				8'b1011001: c <= 9'b111101101;
				8'b110100: c <= 9'b10;
				8'b1111001: c <= 9'b11010100;
				8'b1110001: c <= 9'b100000011;
				8'b1001111: c <= 9'b111100110;
				8'b1100101: c <= 9'b110100100;
				8'b1111110: c <= 9'b11101100;
				8'b1111100: c <= 9'b110000101;
				8'b1010110: c <= 9'b101111110;
				8'b110010: c <= 9'b101;
				8'b1101101: c <= 9'b110100010;
				8'b100011: c <= 9'b11011011;
				8'b1110101: c <= 9'b10100100;
				8'b1111101: c <= 9'b1101110;
				8'b101001: c <= 9'b10000001;
				8'b1010010: c <= 9'b101101100;
				8'b1011000: c <= 9'b110100000;
				8'b101110: c <= 9'b11110101;
				8'b1000001: c <= 9'b111111110;
				default: c <= 9'b0;
			endcase
			9'b101001100 : case(di)
				8'b1000011: c <= 9'b111001011;
				8'b101000: c <= 9'b11;
				8'b111010: c <= 9'b10011000;
				8'b110110: c <= 9'b111000101;
				8'b1100100: c <= 9'b101010000;
				8'b1000000: c <= 9'b100011000;
				8'b1110110: c <= 9'b11110001;
				8'b100101: c <= 9'b111101;
				8'b101111: c <= 9'b11011100;
				8'b100110: c <= 9'b11000100;
				8'b1100011: c <= 9'b10010100;
				8'b1001000: c <= 9'b1011001;
				8'b111000: c <= 9'b101110111;
				8'b110001: c <= 9'b1111101;
				8'b1010111: c <= 9'b111111101;
				8'b1001110: c <= 9'b100000100;
				8'b1101010: c <= 9'b1011110;
				8'b1001001: c <= 9'b10100000;
				8'b1100000: c <= 9'b110000111;
				8'b110111: c <= 9'b100111000;
				8'b1011101: c <= 9'b11111101;
				8'b1011011: c <= 9'b11;
				8'b111001: c <= 9'b1110101;
				8'b1001010: c <= 9'b11100111;
				8'b110011: c <= 9'b111011;
				8'b1101100: c <= 9'b110111010;
				8'b1110111: c <= 9'b11010000;
				8'b101011: c <= 9'b11010101;
				8'b1101011: c <= 9'b10110101;
				8'b111100: c <= 9'b111010111;
				8'b1000111: c <= 9'b101010111;
				8'b1011111: c <= 9'b101101101;
				8'b1110100: c <= 9'b1111111;
				8'b101101: c <= 9'b10000110;
				8'b1010011: c <= 9'b100111;
				8'b1100001: c <= 9'b111111011;
				8'b110101: c <= 9'b10010000;
				8'b1000100: c <= 9'b100111110;
				8'b1010001: c <= 9'b101100010;
				8'b1010100: c <= 9'b1100000;
				8'b1100110: c <= 9'b111100010;
				8'b101010: c <= 9'b111101110;
				8'b1011110: c <= 9'b1110111;
				8'b1100111: c <= 9'b101000101;
				8'b1011010: c <= 9'b1100001;
				8'b1000010: c <= 9'b111010;
				8'b111101: c <= 9'b111001001;
				8'b110000: c <= 9'b11101;
				8'b111110: c <= 9'b100011001;
				8'b1100010: c <= 9'b101100100;
				8'b1110000: c <= 9'b110110000;
				8'b1101001: c <= 9'b10101;
				8'b1110011: c <= 9'b1010101;
				8'b1001100: c <= 9'b111100010;
				8'b100001: c <= 9'b10101100;
				8'b1000110: c <= 9'b110011;
				8'b1110010: c <= 9'b100011011;
				8'b1010000: c <= 9'b111100100;
				8'b1111010: c <= 9'b110101100;
				8'b1010101: c <= 9'b100111111;
				8'b111011: c <= 9'b100000000;
				8'b1001101: c <= 9'b100101000;
				8'b111111: c <= 9'b1011100;
				8'b1101110: c <= 9'b1001011;
				8'b1111011: c <= 9'b111000011;
				8'b1001011: c <= 9'b1110011;
				8'b1101111: c <= 9'b100001001;
				8'b1101000: c <= 9'b10111110;
				8'b101100: c <= 9'b1000100;
				8'b100100: c <= 9'b100111010;
				8'b1111000: c <= 9'b110010100;
				8'b1000101: c <= 9'b10010110;
				8'b1011001: c <= 9'b111101100;
				8'b110100: c <= 9'b110011110;
				8'b1111001: c <= 9'b111001000;
				8'b1110001: c <= 9'b111101100;
				8'b1001111: c <= 9'b100000101;
				8'b1100101: c <= 9'b101110101;
				8'b1111110: c <= 9'b110010100;
				8'b1111100: c <= 9'b101010;
				8'b1010110: c <= 9'b110110110;
				8'b110010: c <= 9'b11000;
				8'b1101101: c <= 9'b1010001;
				8'b100011: c <= 9'b110100110;
				8'b1110101: c <= 9'b101000001;
				8'b1111101: c <= 9'b10001100;
				8'b101001: c <= 9'b1101110;
				8'b1010010: c <= 9'b111111011;
				8'b1011000: c <= 9'b111001010;
				8'b101110: c <= 9'b100111000;
				8'b1000001: c <= 9'b111000110;
				default: c <= 9'b0;
			endcase
			9'b110001 : case(di)
				8'b1000011: c <= 9'b10010110;
				8'b101000: c <= 9'b101010011;
				8'b111010: c <= 9'b11101100;
				8'b110110: c <= 9'b111110001;
				8'b1100100: c <= 9'b11111010;
				8'b1000000: c <= 9'b100000011;
				8'b1110110: c <= 9'b101110;
				8'b100101: c <= 9'b101101010;
				8'b101111: c <= 9'b110001010;
				8'b100110: c <= 9'b1110;
				8'b1100011: c <= 9'b101110011;
				8'b1001000: c <= 9'b110110110;
				8'b111000: c <= 9'b10110;
				8'b110001: c <= 9'b11101;
				8'b1010111: c <= 9'b110011111;
				8'b1001110: c <= 9'b110000010;
				8'b1101010: c <= 9'b111000000;
				8'b1001001: c <= 9'b100111001;
				8'b1100000: c <= 9'b10001101;
				8'b110111: c <= 9'b111001110;
				8'b1011101: c <= 9'b11101000;
				8'b1011011: c <= 9'b10111;
				8'b111001: c <= 9'b11101100;
				8'b1001010: c <= 9'b110000011;
				8'b110011: c <= 9'b1100110;
				8'b1101100: c <= 9'b100101101;
				8'b1110111: c <= 9'b1001100;
				8'b101011: c <= 9'b100100001;
				8'b1101011: c <= 9'b10101;
				8'b111100: c <= 9'b101011001;
				8'b1000111: c <= 9'b101000;
				8'b1011111: c <= 9'b110010011;
				8'b1110100: c <= 9'b100011010;
				8'b101101: c <= 9'b100000001;
				8'b1010011: c <= 9'b11010000;
				8'b1100001: c <= 9'b101111111;
				8'b110101: c <= 9'b110110010;
				8'b1000100: c <= 9'b10110101;
				8'b1010001: c <= 9'b10010000;
				8'b1010100: c <= 9'b1001000;
				8'b1100110: c <= 9'b101010010;
				8'b101010: c <= 9'b1000001;
				8'b1011110: c <= 9'b1001111;
				8'b1100111: c <= 9'b101110;
				8'b1011010: c <= 9'b100001100;
				8'b1000010: c <= 9'b101001000;
				8'b111101: c <= 9'b101111001;
				8'b110000: c <= 9'b11101101;
				8'b111110: c <= 9'b100011001;
				8'b1100010: c <= 9'b11000001;
				8'b1110000: c <= 9'b101010011;
				8'b1101001: c <= 9'b10110100;
				8'b1110011: c <= 9'b100110110;
				8'b1001100: c <= 9'b111010000;
				8'b100001: c <= 9'b11101111;
				8'b1000110: c <= 9'b1111010;
				8'b1110010: c <= 9'b100110000;
				8'b1010000: c <= 9'b10001100;
				8'b1111010: c <= 9'b11110101;
				8'b1010101: c <= 9'b100101101;
				8'b111011: c <= 9'b100000101;
				8'b1001101: c <= 9'b110011101;
				8'b111111: c <= 9'b100111011;
				8'b1101110: c <= 9'b110110010;
				8'b1111011: c <= 9'b1101000;
				8'b1001011: c <= 9'b101110010;
				8'b1101111: c <= 9'b101110110;
				8'b1101000: c <= 9'b111100110;
				8'b101100: c <= 9'b100100000;
				8'b100100: c <= 9'b11110111;
				8'b1111000: c <= 9'b1;
				8'b1000101: c <= 9'b101101010;
				8'b1011001: c <= 9'b1011110;
				8'b110100: c <= 9'b110110111;
				8'b1111001: c <= 9'b111011010;
				8'b1110001: c <= 9'b101110110;
				8'b1001111: c <= 9'b10110101;
				8'b1100101: c <= 9'b110000111;
				8'b1111110: c <= 9'b110000001;
				8'b1111100: c <= 9'b10010011;
				8'b1010110: c <= 9'b11110010;
				8'b110010: c <= 9'b111100101;
				8'b1101101: c <= 9'b101111000;
				8'b100011: c <= 9'b10010011;
				8'b1110101: c <= 9'b111111011;
				8'b1111101: c <= 9'b100111100;
				8'b101001: c <= 9'b111010001;
				8'b1010010: c <= 9'b111110011;
				8'b1011000: c <= 9'b111011110;
				8'b101110: c <= 9'b1100000;
				8'b1000001: c <= 9'b1000111;
				default: c <= 9'b0;
			endcase
			9'b111011101 : case(di)
				8'b1000011: c <= 9'b110011010;
				8'b101000: c <= 9'b1001101;
				8'b111010: c <= 9'b111000010;
				8'b110110: c <= 9'b11001111;
				8'b1100100: c <= 9'b1000000;
				8'b1000000: c <= 9'b111110110;
				8'b1110110: c <= 9'b100111110;
				8'b100101: c <= 9'b110100000;
				8'b101111: c <= 9'b1001010;
				8'b100110: c <= 9'b1000011;
				8'b1100011: c <= 9'b100010100;
				8'b1001000: c <= 9'b10101000;
				8'b111000: c <= 9'b111100110;
				8'b110001: c <= 9'b11000110;
				8'b1010111: c <= 9'b100111001;
				8'b1001110: c <= 9'b1110;
				8'b1101010: c <= 9'b11001111;
				8'b1001001: c <= 9'b11110111;
				8'b1100000: c <= 9'b11010011;
				8'b110111: c <= 9'b111110000;
				8'b1011101: c <= 9'b100000011;
				8'b1011011: c <= 9'b100100010;
				8'b111001: c <= 9'b110101110;
				8'b1001010: c <= 9'b1010010;
				8'b110011: c <= 9'b100110;
				8'b1101100: c <= 9'b11101100;
				8'b1110111: c <= 9'b111101001;
				8'b101011: c <= 9'b10010101;
				8'b1101011: c <= 9'b110001111;
				8'b111100: c <= 9'b101110100;
				8'b1000111: c <= 9'b10;
				8'b1011111: c <= 9'b101111111;
				8'b1110100: c <= 9'b111100000;
				8'b101101: c <= 9'b11001001;
				8'b1010011: c <= 9'b110100110;
				8'b1100001: c <= 9'b111000011;
				8'b110101: c <= 9'b111011;
				8'b1000100: c <= 9'b1110010;
				8'b1010001: c <= 9'b100101101;
				8'b1010100: c <= 9'b10101;
				8'b1100110: c <= 9'b110110111;
				8'b101010: c <= 9'b110110;
				8'b1011110: c <= 9'b1010011;
				8'b1100111: c <= 9'b101000101;
				8'b1011010: c <= 9'b101010100;
				8'b1000010: c <= 9'b11011101;
				8'b111101: c <= 9'b100001111;
				8'b110000: c <= 9'b10100011;
				8'b111110: c <= 9'b11010;
				8'b1100010: c <= 9'b1010101;
				8'b1110000: c <= 9'b111101000;
				8'b1101001: c <= 9'b10110;
				8'b1110011: c <= 9'b101010100;
				8'b1001100: c <= 9'b11110000;
				8'b100001: c <= 9'b111001100;
				8'b1000110: c <= 9'b101010111;
				8'b1110010: c <= 9'b110101010;
				8'b1010000: c <= 9'b111010110;
				8'b1111010: c <= 9'b1000111;
				8'b1010101: c <= 9'b101010110;
				8'b111011: c <= 9'b1110000;
				8'b1001101: c <= 9'b10001110;
				8'b111111: c <= 9'b10100100;
				8'b1101110: c <= 9'b10000000;
				8'b1111011: c <= 9'b11110100;
				8'b1001011: c <= 9'b111000011;
				8'b1101111: c <= 9'b100111000;
				8'b1101000: c <= 9'b11110100;
				8'b101100: c <= 9'b10111100;
				8'b100100: c <= 9'b111001001;
				8'b1111000: c <= 9'b101100100;
				8'b1000101: c <= 9'b110111;
				8'b1011001: c <= 9'b1111110;
				8'b110100: c <= 9'b101101;
				8'b1111001: c <= 9'b11111001;
				8'b1110001: c <= 9'b110011011;
				8'b1001111: c <= 9'b10110010;
				8'b1100101: c <= 9'b100110110;
				8'b1111110: c <= 9'b110000011;
				8'b1111100: c <= 9'b11111001;
				8'b1010110: c <= 9'b111011011;
				8'b110010: c <= 9'b10011;
				8'b1101101: c <= 9'b111010110;
				8'b100011: c <= 9'b1;
				8'b1110101: c <= 9'b111000110;
				8'b1111101: c <= 9'b101101011;
				8'b101001: c <= 9'b1001110;
				8'b1010010: c <= 9'b1011010;
				8'b1011000: c <= 9'b10110;
				8'b101110: c <= 9'b111101101;
				8'b1000001: c <= 9'b10001111;
				default: c <= 9'b0;
			endcase
			9'b11100101 : case(di)
				8'b1000011: c <= 9'b10111;
				8'b101000: c <= 9'b111001110;
				8'b111010: c <= 9'b111000010;
				8'b110110: c <= 9'b100111011;
				8'b1100100: c <= 9'b110010010;
				8'b1000000: c <= 9'b1000;
				8'b1110110: c <= 9'b110010101;
				8'b100101: c <= 9'b110100111;
				8'b101111: c <= 9'b101010111;
				8'b100110: c <= 9'b100111110;
				8'b1100011: c <= 9'b111101101;
				8'b1001000: c <= 9'b1101111;
				8'b111000: c <= 9'b11011101;
				8'b110001: c <= 9'b110100101;
				8'b1010111: c <= 9'b100111110;
				8'b1001110: c <= 9'b10000101;
				8'b1101010: c <= 9'b110000001;
				8'b1001001: c <= 9'b10011010;
				8'b1100000: c <= 9'b10000011;
				8'b110111: c <= 9'b10001010;
				8'b1011101: c <= 9'b100100111;
				8'b1011011: c <= 9'b100010100;
				8'b111001: c <= 9'b110011010;
				8'b1001010: c <= 9'b111000000;
				8'b110011: c <= 9'b11110110;
				8'b1101100: c <= 9'b111111110;
				8'b1110111: c <= 9'b111001010;
				8'b101011: c <= 9'b10110001;
				8'b1101011: c <= 9'b10001010;
				8'b111100: c <= 9'b111100010;
				8'b1000111: c <= 9'b101110010;
				8'b1011111: c <= 9'b1010111;
				8'b1110100: c <= 9'b110001010;
				8'b101101: c <= 9'b101;
				8'b1010011: c <= 9'b110001011;
				8'b1100001: c <= 9'b1011;
				8'b110101: c <= 9'b100000010;
				8'b1000100: c <= 9'b11110000;
				8'b1010001: c <= 9'b10110011;
				8'b1010100: c <= 9'b101100;
				8'b1100110: c <= 9'b101010;
				8'b101010: c <= 9'b100111;
				8'b1011110: c <= 9'b111101000;
				8'b1100111: c <= 9'b111001110;
				8'b1011010: c <= 9'b1010111;
				8'b1000010: c <= 9'b1001000;
				8'b111101: c <= 9'b11100100;
				8'b110000: c <= 9'b10010110;
				8'b111110: c <= 9'b100010110;
				8'b1100010: c <= 9'b1101101;
				8'b1110000: c <= 9'b110110;
				8'b1101001: c <= 9'b100001111;
				8'b1110011: c <= 9'b111001101;
				8'b1001100: c <= 9'b110100001;
				8'b100001: c <= 9'b110000111;
				8'b1000110: c <= 9'b11000010;
				8'b1110010: c <= 9'b11111110;
				8'b1010000: c <= 9'b100111000;
				8'b1111010: c <= 9'b110101101;
				8'b1010101: c <= 9'b101100111;
				8'b111011: c <= 9'b110011000;
				8'b1001101: c <= 9'b101000110;
				8'b111111: c <= 9'b10011100;
				8'b1101110: c <= 9'b110110101;
				8'b1111011: c <= 9'b111011110;
				8'b1001011: c <= 9'b111111001;
				8'b1101111: c <= 9'b11011010;
				8'b1101000: c <= 9'b1010111;
				8'b101100: c <= 9'b111000101;
				8'b100100: c <= 9'b10001111;
				8'b1111000: c <= 9'b110010010;
				8'b1000101: c <= 9'b111101101;
				8'b1011001: c <= 9'b10001011;
				8'b110100: c <= 9'b110101011;
				8'b1111001: c <= 9'b100111010;
				8'b1110001: c <= 9'b101101001;
				8'b1001111: c <= 9'b11001001;
				8'b1100101: c <= 9'b110000110;
				8'b1111110: c <= 9'b110011101;
				8'b1111100: c <= 9'b100101100;
				8'b1010110: c <= 9'b101111001;
				8'b110010: c <= 9'b10011100;
				8'b1101101: c <= 9'b101000001;
				8'b100011: c <= 9'b101110111;
				8'b1110101: c <= 9'b100011011;
				8'b1111101: c <= 9'b10101011;
				8'b101001: c <= 9'b110101011;
				8'b1010010: c <= 9'b110011111;
				8'b1011000: c <= 9'b10;
				8'b101110: c <= 9'b111000100;
				8'b1000001: c <= 9'b100010111;
				default: c <= 9'b0;
			endcase
			9'b10100000 : case(di)
				8'b1000011: c <= 9'b100101010;
				8'b101000: c <= 9'b110010010;
				8'b111010: c <= 9'b111000;
				8'b110110: c <= 9'b100000011;
				8'b1100100: c <= 9'b1000010;
				8'b1000000: c <= 9'b101010000;
				8'b1110110: c <= 9'b100101011;
				8'b100101: c <= 9'b101001000;
				8'b101111: c <= 9'b10111101;
				8'b100110: c <= 9'b100100110;
				8'b1100011: c <= 9'b101011101;
				8'b1001000: c <= 9'b101010010;
				8'b111000: c <= 9'b10001100;
				8'b110001: c <= 9'b10011001;
				8'b1010111: c <= 9'b1001100;
				8'b1001110: c <= 9'b11110000;
				8'b1101010: c <= 9'b10001100;
				8'b1001001: c <= 9'b110111110;
				8'b1100000: c <= 9'b111011001;
				8'b110111: c <= 9'b100011000;
				8'b1011101: c <= 9'b1110100;
				8'b1011011: c <= 9'b111110011;
				8'b111001: c <= 9'b10100110;
				8'b1001010: c <= 9'b10000111;
				8'b110011: c <= 9'b110110100;
				8'b1101100: c <= 9'b11011010;
				8'b1110111: c <= 9'b110001011;
				8'b101011: c <= 9'b111101101;
				8'b1101011: c <= 9'b11010001;
				8'b111100: c <= 9'b111;
				8'b1000111: c <= 9'b11100010;
				8'b1011111: c <= 9'b11011;
				8'b1110100: c <= 9'b1101111;
				8'b101101: c <= 9'b100100101;
				8'b1010011: c <= 9'b111011110;
				8'b1100001: c <= 9'b110010011;
				8'b110101: c <= 9'b101100010;
				8'b1000100: c <= 9'b100111001;
				8'b1010001: c <= 9'b11001;
				8'b1010100: c <= 9'b1000010;
				8'b1100110: c <= 9'b101111111;
				8'b101010: c <= 9'b100001010;
				8'b1011110: c <= 9'b101011110;
				8'b1100111: c <= 9'b10100111;
				8'b1011010: c <= 9'b100000111;
				8'b1000010: c <= 9'b1100111;
				8'b111101: c <= 9'b110101110;
				8'b110000: c <= 9'b10000001;
				8'b111110: c <= 9'b111000;
				8'b1100010: c <= 9'b110101001;
				8'b1110000: c <= 9'b1110000;
				8'b1101001: c <= 9'b10111000;
				8'b1110011: c <= 9'b11011000;
				8'b1001100: c <= 9'b100100111;
				8'b100001: c <= 9'b100011101;
				8'b1000110: c <= 9'b11010000;
				8'b1110010: c <= 9'b1101001;
				8'b1010000: c <= 9'b11011011;
				8'b1111010: c <= 9'b11011;
				8'b1010101: c <= 9'b111011010;
				8'b111011: c <= 9'b1111101;
				8'b1001101: c <= 9'b10100111;
				8'b111111: c <= 9'b110101011;
				8'b1101110: c <= 9'b110110010;
				8'b1111011: c <= 9'b111000000;
				8'b1001011: c <= 9'b100101001;
				8'b1101111: c <= 9'b110111010;
				8'b1101000: c <= 9'b10111010;
				8'b101100: c <= 9'b111001010;
				8'b100100: c <= 9'b101101101;
				8'b1111000: c <= 9'b110100001;
				8'b1000101: c <= 9'b111000111;
				8'b1011001: c <= 9'b110111100;
				8'b110100: c <= 9'b111000010;
				8'b1111001: c <= 9'b111010001;
				8'b1110001: c <= 9'b101100010;
				8'b1001111: c <= 9'b111111000;
				8'b1100101: c <= 9'b101101010;
				8'b1111110: c <= 9'b101000011;
				8'b1111100: c <= 9'b1111010;
				8'b1010110: c <= 9'b11100011;
				8'b110010: c <= 9'b101111001;
				8'b1101101: c <= 9'b110011000;
				8'b100011: c <= 9'b111100;
				8'b1110101: c <= 9'b111011101;
				8'b1111101: c <= 9'b111001001;
				8'b101001: c <= 9'b101110000;
				8'b1010010: c <= 9'b1111000;
				8'b1011000: c <= 9'b11010100;
				8'b101110: c <= 9'b1100101;
				8'b1000001: c <= 9'b100000101;
				default: c <= 9'b0;
			endcase
			9'b111001 : case(di)
				8'b1000011: c <= 9'b111111000;
				8'b101000: c <= 9'b111101;
				8'b111010: c <= 9'b111;
				8'b110110: c <= 9'b100101010;
				8'b1100100: c <= 9'b11001101;
				8'b1000000: c <= 9'b110001001;
				8'b1110110: c <= 9'b111100111;
				8'b100101: c <= 9'b11000110;
				8'b101111: c <= 9'b100000110;
				8'b100110: c <= 9'b110011100;
				8'b1100011: c <= 9'b111110001;
				8'b1001000: c <= 9'b100111100;
				8'b111000: c <= 9'b100111101;
				8'b110001: c <= 9'b1000000;
				8'b1010111: c <= 9'b10000000;
				8'b1001110: c <= 9'b10001010;
				8'b1101010: c <= 9'b1100010;
				8'b1001001: c <= 9'b100101;
				8'b1100000: c <= 9'b100011001;
				8'b110111: c <= 9'b1110111;
				8'b1011101: c <= 9'b111000011;
				8'b1011011: c <= 9'b111000011;
				8'b111001: c <= 9'b10000110;
				8'b1001010: c <= 9'b100011010;
				8'b110011: c <= 9'b100001100;
				8'b1101100: c <= 9'b10101000;
				8'b1110111: c <= 9'b1001110;
				8'b101011: c <= 9'b11110111;
				8'b1101011: c <= 9'b11100110;
				8'b111100: c <= 9'b100011101;
				8'b1000111: c <= 9'b100000000;
				8'b1011111: c <= 9'b1110111;
				8'b1110100: c <= 9'b100101001;
				8'b101101: c <= 9'b101011010;
				8'b1010011: c <= 9'b1110;
				8'b1100001: c <= 9'b101111001;
				8'b110101: c <= 9'b100101101;
				8'b1000100: c <= 9'b10001100;
				8'b1010001: c <= 9'b110000000;
				8'b1010100: c <= 9'b10000000;
				8'b1100110: c <= 9'b110101100;
				8'b101010: c <= 9'b101000011;
				8'b1011110: c <= 9'b110000010;
				8'b1100111: c <= 9'b11101011;
				8'b1011010: c <= 9'b1010000;
				8'b1000010: c <= 9'b11001100;
				8'b111101: c <= 9'b101010011;
				8'b110000: c <= 9'b1110000;
				8'b111110: c <= 9'b10111000;
				8'b1100010: c <= 9'b10111011;
				8'b1110000: c <= 9'b10101110;
				8'b1101001: c <= 9'b101001;
				8'b1110011: c <= 9'b10101100;
				8'b1001100: c <= 9'b100111100;
				8'b100001: c <= 9'b1000110;
				8'b1000110: c <= 9'b10111110;
				8'b1110010: c <= 9'b11000;
				8'b1010000: c <= 9'b101100011;
				8'b1111010: c <= 9'b10100111;
				8'b1010101: c <= 9'b1001110;
				8'b111011: c <= 9'b100100101;
				8'b1001101: c <= 9'b11110;
				8'b111111: c <= 9'b10011001;
				8'b1101110: c <= 9'b101111110;
				8'b1111011: c <= 9'b111101100;
				8'b1001011: c <= 9'b110111011;
				8'b1101111: c <= 9'b110100010;
				8'b1101000: c <= 9'b110100010;
				8'b101100: c <= 9'b100110;
				8'b100100: c <= 9'b1010001;
				8'b1111000: c <= 9'b1110000;
				8'b1000101: c <= 9'b111001111;
				8'b1011001: c <= 9'b101011010;
				8'b110100: c <= 9'b100001110;
				8'b1111001: c <= 9'b110110;
				8'b1110001: c <= 9'b10010000;
				8'b1001111: c <= 9'b100101111;
				8'b1100101: c <= 9'b1010000;
				8'b1111110: c <= 9'b11;
				8'b1111100: c <= 9'b110011;
				8'b1010110: c <= 9'b1011;
				8'b110010: c <= 9'b1000111;
				8'b1101101: c <= 9'b11010001;
				8'b100011: c <= 9'b101000110;
				8'b1110101: c <= 9'b11010;
				8'b1111101: c <= 9'b1100;
				8'b101001: c <= 9'b1001111;
				8'b1010010: c <= 9'b111001110;
				8'b1011000: c <= 9'b101100101;
				8'b101110: c <= 9'b100001110;
				8'b1000001: c <= 9'b111001110;
				default: c <= 9'b0;
			endcase
			9'b1111100 : case(di)
				8'b1000011: c <= 9'b110010110;
				8'b101000: c <= 9'b10011101;
				8'b111010: c <= 9'b101001001;
				8'b110110: c <= 9'b100101;
				8'b1100100: c <= 9'b1100001;
				8'b1000000: c <= 9'b101101;
				8'b1110110: c <= 9'b111010;
				8'b100101: c <= 9'b1110011;
				8'b101111: c <= 9'b111011101;
				8'b100110: c <= 9'b11011100;
				8'b1100011: c <= 9'b11101100;
				8'b1001000: c <= 9'b10101110;
				8'b111000: c <= 9'b11000000;
				8'b110001: c <= 9'b101001;
				8'b1010111: c <= 9'b1010101;
				8'b1001110: c <= 9'b101110111;
				8'b1101010: c <= 9'b10001100;
				8'b1001001: c <= 9'b110000111;
				8'b1100000: c <= 9'b110000001;
				8'b110111: c <= 9'b11110000;
				8'b1011101: c <= 9'b101100110;
				8'b1011011: c <= 9'b110110101;
				8'b111001: c <= 9'b11000000;
				8'b1001010: c <= 9'b110010100;
				8'b110011: c <= 9'b11011110;
				8'b1101100: c <= 9'b11111011;
				8'b1110111: c <= 9'b100010101;
				8'b101011: c <= 9'b100011000;
				8'b1101011: c <= 9'b110100100;
				8'b111100: c <= 9'b101101110;
				8'b1000111: c <= 9'b111110101;
				8'b1011111: c <= 9'b1010000;
				8'b1110100: c <= 9'b100100110;
				8'b101101: c <= 9'b101111110;
				8'b1010011: c <= 9'b11110110;
				8'b1100001: c <= 9'b100111;
				8'b110101: c <= 9'b10010111;
				8'b1000100: c <= 9'b10000110;
				8'b1010001: c <= 9'b101100111;
				8'b1010100: c <= 9'b1010010;
				8'b1100110: c <= 9'b110011110;
				8'b101010: c <= 9'b11001100;
				8'b1011110: c <= 9'b11011101;
				8'b1100111: c <= 9'b11000001;
				8'b1011010: c <= 9'b111111101;
				8'b1000010: c <= 9'b10001010;
				8'b111101: c <= 9'b10010;
				8'b110000: c <= 9'b11010101;
				8'b111110: c <= 9'b111100101;
				8'b1100010: c <= 9'b110010001;
				8'b1110000: c <= 9'b11101011;
				8'b1101001: c <= 9'b111101001;
				8'b1110011: c <= 9'b101100101;
				8'b1001100: c <= 9'b10100000;
				8'b100001: c <= 9'b1010111;
				8'b1000110: c <= 9'b100101000;
				8'b1110010: c <= 9'b111010010;
				8'b1010000: c <= 9'b1011110;
				8'b1111010: c <= 9'b110100;
				8'b1010101: c <= 9'b1101001;
				8'b111011: c <= 9'b1111001;
				8'b1001101: c <= 9'b110101001;
				8'b111111: c <= 9'b110010001;
				8'b1101110: c <= 9'b101100011;
				8'b1111011: c <= 9'b101011111;
				8'b1001011: c <= 9'b10001100;
				8'b1101111: c <= 9'b1110000;
				8'b1101000: c <= 9'b1010010;
				8'b101100: c <= 9'b1001001;
				8'b100100: c <= 9'b101111110;
				8'b1111000: c <= 9'b10011010;
				8'b1000101: c <= 9'b101110111;
				8'b1011001: c <= 9'b110001100;
				8'b110100: c <= 9'b10001001;
				8'b1111001: c <= 9'b11110;
				8'b1110001: c <= 9'b1100010;
				8'b1001111: c <= 9'b101010111;
				8'b1100101: c <= 9'b100110100;
				8'b1111110: c <= 9'b100111011;
				8'b1111100: c <= 9'b111111001;
				8'b1010110: c <= 9'b100110011;
				8'b110010: c <= 9'b100010100;
				8'b1101101: c <= 9'b110010011;
				8'b100011: c <= 9'b1011100;
				8'b1110101: c <= 9'b1100001;
				8'b1111101: c <= 9'b11101011;
				8'b101001: c <= 9'b10011011;
				8'b1010010: c <= 9'b101101;
				8'b1011000: c <= 9'b10011010;
				8'b101110: c <= 9'b110011010;
				8'b1000001: c <= 9'b111100011;
				default: c <= 9'b0;
			endcase
			9'b10 : case(di)
				8'b1000011: c <= 9'b110001101;
				8'b101000: c <= 9'b10000000;
				8'b111010: c <= 9'b111011111;
				8'b110110: c <= 9'b111001111;
				8'b1100100: c <= 9'b110010;
				8'b1000000: c <= 9'b11001101;
				8'b1110110: c <= 9'b1100;
				8'b100101: c <= 9'b110011010;
				8'b101111: c <= 9'b1110010;
				8'b100110: c <= 9'b100011;
				8'b1100011: c <= 9'b110111010;
				8'b1001000: c <= 9'b111111110;
				8'b111000: c <= 9'b101001;
				8'b110001: c <= 9'b11110111;
				8'b1010111: c <= 9'b101101010;
				8'b1001110: c <= 9'b111101000;
				8'b1101010: c <= 9'b100101100;
				8'b1001001: c <= 9'b101010111;
				8'b1100000: c <= 9'b10011;
				8'b110111: c <= 9'b1111111;
				8'b1011101: c <= 9'b100011101;
				8'b1011011: c <= 9'b1000011;
				8'b111001: c <= 9'b11010000;
				8'b1001010: c <= 9'b1011;
				8'b110011: c <= 9'b110100000;
				8'b1101100: c <= 9'b100101011;
				8'b1110111: c <= 9'b1101100;
				8'b101011: c <= 9'b111;
				8'b1101011: c <= 9'b1111101;
				8'b111100: c <= 9'b11001011;
				8'b1000111: c <= 9'b111000111;
				8'b1011111: c <= 9'b11000111;
				8'b1110100: c <= 9'b100011101;
				8'b101101: c <= 9'b100110111;
				8'b1010011: c <= 9'b110110011;
				8'b1100001: c <= 9'b110101001;
				8'b110101: c <= 9'b110110100;
				8'b1000100: c <= 9'b111100100;
				8'b1010001: c <= 9'b1011001;
				8'b1010100: c <= 9'b110011000;
				8'b1100110: c <= 9'b11111;
				8'b101010: c <= 9'b1001011;
				8'b1011110: c <= 9'b11010000;
				8'b1100111: c <= 9'b11101;
				8'b1011010: c <= 9'b1101010;
				8'b1000010: c <= 9'b10110011;
				8'b111101: c <= 9'b101100100;
				8'b110000: c <= 9'b10010;
				8'b111110: c <= 9'b111010001;
				8'b1100010: c <= 9'b111001101;
				8'b1110000: c <= 9'b101110100;
				8'b1101001: c <= 9'b1111000;
				8'b1110011: c <= 9'b10111100;
				8'b1001100: c <= 9'b1010101;
				8'b100001: c <= 9'b110101;
				8'b1000110: c <= 9'b10000110;
				8'b1110010: c <= 9'b1011111;
				8'b1010000: c <= 9'b111001000;
				8'b1111010: c <= 9'b1001100;
				8'b1010101: c <= 9'b1101001;
				8'b111011: c <= 9'b111110000;
				8'b1001101: c <= 9'b10110111;
				8'b111111: c <= 9'b111001101;
				8'b1101110: c <= 9'b110000000;
				8'b1111011: c <= 9'b10000011;
				8'b1001011: c <= 9'b11001100;
				8'b1101111: c <= 9'b11001010;
				8'b1101000: c <= 9'b11001010;
				8'b101100: c <= 9'b101100111;
				8'b100100: c <= 9'b100100111;
				8'b1111000: c <= 9'b1110;
				8'b1000101: c <= 9'b100101000;
				8'b1011001: c <= 9'b111011101;
				8'b110100: c <= 9'b100101101;
				8'b1111001: c <= 9'b100000110;
				8'b1110001: c <= 9'b110010;
				8'b1001111: c <= 9'b100100101;
				8'b1100101: c <= 9'b101111010;
				8'b1111110: c <= 9'b101111110;
				8'b1111100: c <= 9'b110011101;
				8'b1010110: c <= 9'b100100001;
				8'b110010: c <= 9'b100011011;
				8'b1101101: c <= 9'b11000001;
				8'b100011: c <= 9'b111110110;
				8'b1110101: c <= 9'b10011011;
				8'b1111101: c <= 9'b100101100;
				8'b101001: c <= 9'b1100110;
				8'b1010010: c <= 9'b10000011;
				8'b1011000: c <= 9'b11010010;
				8'b101110: c <= 9'b10001000;
				8'b1000001: c <= 9'b110;
				default: c <= 9'b0;
			endcase
			9'b111110011 : case(di)
				8'b1000011: c <= 9'b101101;
				8'b101000: c <= 9'b10110110;
				8'b111010: c <= 9'b100110010;
				8'b110110: c <= 9'b100111001;
				8'b1100100: c <= 9'b111111;
				8'b1000000: c <= 9'b11001011;
				8'b1110110: c <= 9'b1111101;
				8'b100101: c <= 9'b1101100;
				8'b101111: c <= 9'b1100001;
				8'b100110: c <= 9'b101011111;
				8'b1100011: c <= 9'b111110000;
				8'b1001000: c <= 9'b101000101;
				8'b111000: c <= 9'b11101000;
				8'b110001: c <= 9'b10100011;
				8'b1010111: c <= 9'b100001011;
				8'b1001110: c <= 9'b11011001;
				8'b1101010: c <= 9'b111110110;
				8'b1001001: c <= 9'b11011011;
				8'b1100000: c <= 9'b1110101;
				8'b110111: c <= 9'b100101100;
				8'b1011101: c <= 9'b110010111;
				8'b1011011: c <= 9'b11001100;
				8'b111001: c <= 9'b10010100;
				8'b1001010: c <= 9'b111100001;
				8'b110011: c <= 9'b111111111;
				8'b1101100: c <= 9'b11100100;
				8'b1110111: c <= 9'b111011011;
				8'b101011: c <= 9'b11010001;
				8'b1101011: c <= 9'b111111010;
				8'b111100: c <= 9'b110011110;
				8'b1000111: c <= 9'b111101110;
				8'b1011111: c <= 9'b10001001;
				8'b1110100: c <= 9'b10010011;
				8'b101101: c <= 9'b11000100;
				8'b1010011: c <= 9'b100110110;
				8'b1100001: c <= 9'b11111011;
				8'b110101: c <= 9'b110011010;
				8'b1000100: c <= 9'b110;
				8'b1010001: c <= 9'b10111110;
				8'b1010100: c <= 9'b111011111;
				8'b1100110: c <= 9'b1111;
				8'b101010: c <= 9'b1011100;
				8'b1011110: c <= 9'b111010000;
				8'b1100111: c <= 9'b111010;
				8'b1011010: c <= 9'b100101101;
				8'b1000010: c <= 9'b1100000;
				8'b111101: c <= 9'b111101010;
				8'b110000: c <= 9'b100101000;
				8'b111110: c <= 9'b111001011;
				8'b1100010: c <= 9'b100101110;
				8'b1110000: c <= 9'b1001001;
				8'b1101001: c <= 9'b10100011;
				8'b1110011: c <= 9'b111001011;
				8'b1001100: c <= 9'b11111101;
				8'b100001: c <= 9'b111100001;
				8'b1000110: c <= 9'b110000001;
				8'b1110010: c <= 9'b110111111;
				8'b1010000: c <= 9'b101010101;
				8'b1111010: c <= 9'b100010111;
				8'b1010101: c <= 9'b10100010;
				8'b111011: c <= 9'b100000001;
				8'b1001101: c <= 9'b1110001;
				8'b111111: c <= 9'b100001101;
				8'b1101110: c <= 9'b100111111;
				8'b1111011: c <= 9'b11001111;
				8'b1001011: c <= 9'b100110110;
				8'b1101111: c <= 9'b1010011;
				8'b1101000: c <= 9'b111011101;
				8'b101100: c <= 9'b1100010;
				8'b100100: c <= 9'b10010;
				8'b1111000: c <= 9'b1101100;
				8'b1000101: c <= 9'b110101011;
				8'b1011001: c <= 9'b101000010;
				8'b110100: c <= 9'b1000101;
				8'b1111001: c <= 9'b10011100;
				8'b1110001: c <= 9'b101111010;
				8'b1001111: c <= 9'b11101101;
				8'b1100101: c <= 9'b100010;
				8'b1111110: c <= 9'b10110101;
				8'b1111100: c <= 9'b10100101;
				8'b1010110: c <= 9'b101001110;
				8'b110010: c <= 9'b101100101;
				8'b1101101: c <= 9'b1011;
				8'b100011: c <= 9'b101101101;
				8'b1110101: c <= 9'b1111001;
				8'b1111101: c <= 9'b111011001;
				8'b101001: c <= 9'b1010101;
				8'b1010010: c <= 9'b1011000;
				8'b1011000: c <= 9'b101001111;
				8'b101110: c <= 9'b11100001;
				8'b1000001: c <= 9'b101001000;
				default: c <= 9'b0;
			endcase
			9'b111010100 : case(di)
				8'b1000011: c <= 9'b10011100;
				8'b101000: c <= 9'b111001;
				8'b111010: c <= 9'b11011010;
				8'b110110: c <= 9'b110001110;
				8'b1100100: c <= 9'b100110010;
				8'b1000000: c <= 9'b100101101;
				8'b1110110: c <= 9'b110101100;
				8'b100101: c <= 9'b11011110;
				8'b101111: c <= 9'b100111100;
				8'b100110: c <= 9'b11111100;
				8'b1100011: c <= 9'b10101000;
				8'b1001000: c <= 9'b111001000;
				8'b111000: c <= 9'b110011101;
				8'b110001: c <= 9'b111110011;
				8'b1010111: c <= 9'b111011010;
				8'b1001110: c <= 9'b10011010;
				8'b1101010: c <= 9'b101000100;
				8'b1001001: c <= 9'b11001100;
				8'b1100000: c <= 9'b11010001;
				8'b110111: c <= 9'b10000011;
				8'b1011101: c <= 9'b1000001;
				8'b1011011: c <= 9'b11001010;
				8'b111001: c <= 9'b1000011;
				8'b1001010: c <= 9'b11101100;
				8'b110011: c <= 9'b10100101;
				8'b1101100: c <= 9'b110111110;
				8'b1110111: c <= 9'b100001;
				8'b101011: c <= 9'b100000000;
				8'b1101011: c <= 9'b110010010;
				8'b111100: c <= 9'b101000101;
				8'b1000111: c <= 9'b11010111;
				8'b1011111: c <= 9'b101101110;
				8'b1110100: c <= 9'b100110000;
				8'b101101: c <= 9'b11011101;
				8'b1010011: c <= 9'b1011100;
				8'b1100001: c <= 9'b111111010;
				8'b110101: c <= 9'b110101010;
				8'b1000100: c <= 9'b1000011;
				8'b1010001: c <= 9'b11010000;
				8'b1010100: c <= 9'b1011;
				8'b1100110: c <= 9'b111101010;
				8'b101010: c <= 9'b1110001;
				8'b1011110: c <= 9'b100101;
				8'b1100111: c <= 9'b10101100;
				8'b1011010: c <= 9'b1100010;
				8'b1000010: c <= 9'b10101111;
				8'b111101: c <= 9'b111101010;
				8'b110000: c <= 9'b10110110;
				8'b111110: c <= 9'b11100000;
				8'b1100010: c <= 9'b111011110;
				8'b1110000: c <= 9'b110011101;
				8'b1101001: c <= 9'b111100011;
				8'b1110011: c <= 9'b1011001;
				8'b1001100: c <= 9'b111000000;
				8'b100001: c <= 9'b11110011;
				8'b1000110: c <= 9'b100110000;
				8'b1110010: c <= 9'b1010110;
				8'b1010000: c <= 9'b111111001;
				8'b1111010: c <= 9'b1011000;
				8'b1010101: c <= 9'b10011010;
				8'b111011: c <= 9'b10110001;
				8'b1001101: c <= 9'b11111;
				8'b111111: c <= 9'b110100011;
				8'b1101110: c <= 9'b11111011;
				8'b1111011: c <= 9'b111101010;
				8'b1001011: c <= 9'b100010111;
				8'b1101111: c <= 9'b11010010;
				8'b1101000: c <= 9'b1001000;
				8'b101100: c <= 9'b1011010;
				8'b100100: c <= 9'b10101110;
				8'b1111000: c <= 9'b1100001;
				8'b1000101: c <= 9'b111000;
				8'b1011001: c <= 9'b101001100;
				8'b110100: c <= 9'b101110000;
				8'b1111001: c <= 9'b11100;
				8'b1110001: c <= 9'b111011010;
				8'b1001111: c <= 9'b100101011;
				8'b1100101: c <= 9'b110010011;
				8'b1111110: c <= 9'b10101010;
				8'b1111100: c <= 9'b110000111;
				8'b1010110: c <= 9'b101001111;
				8'b110010: c <= 9'b10000000;
				8'b1101101: c <= 9'b100110011;
				8'b100011: c <= 9'b10110010;
				8'b1110101: c <= 9'b101101101;
				8'b1111101: c <= 9'b100100000;
				8'b101001: c <= 9'b1000001;
				8'b1010010: c <= 9'b1110101;
				8'b1011000: c <= 9'b1001111;
				8'b101110: c <= 9'b1101010;
				8'b1000001: c <= 9'b11111110;
				default: c <= 9'b0;
			endcase
			9'b100110000 : case(di)
				8'b1000011: c <= 9'b11111;
				8'b101000: c <= 9'b110000011;
				8'b111010: c <= 9'b101000100;
				8'b110110: c <= 9'b110001000;
				8'b1100100: c <= 9'b111;
				8'b1000000: c <= 9'b100100110;
				8'b1110110: c <= 9'b100111100;
				8'b100101: c <= 9'b11110111;
				8'b101111: c <= 9'b11011100;
				8'b100110: c <= 9'b1100010;
				8'b1100011: c <= 9'b11010101;
				8'b1001000: c <= 9'b110010010;
				8'b111000: c <= 9'b10100111;
				8'b110001: c <= 9'b100101110;
				8'b1010111: c <= 9'b101010111;
				8'b1001110: c <= 9'b101110001;
				8'b1101010: c <= 9'b111001;
				8'b1001001: c <= 9'b111111010;
				8'b1100000: c <= 9'b110100001;
				8'b110111: c <= 9'b100101110;
				8'b1011101: c <= 9'b10010110;
				8'b1011011: c <= 9'b11001011;
				8'b111001: c <= 9'b100100010;
				8'b1001010: c <= 9'b110000110;
				8'b110011: c <= 9'b110101101;
				8'b1101100: c <= 9'b1010001;
				8'b1110111: c <= 9'b11011010;
				8'b101011: c <= 9'b110111011;
				8'b1101011: c <= 9'b110010011;
				8'b111100: c <= 9'b11101;
				8'b1000111: c <= 9'b10000111;
				8'b1011111: c <= 9'b110000111;
				8'b1110100: c <= 9'b10111000;
				8'b101101: c <= 9'b101000001;
				8'b1010011: c <= 9'b100001011;
				8'b1100001: c <= 9'b1111110;
				8'b110101: c <= 9'b10000000;
				8'b1000100: c <= 9'b10001011;
				8'b1010001: c <= 9'b1100001;
				8'b1010100: c <= 9'b1110011;
				8'b1100110: c <= 9'b111110011;
				8'b101010: c <= 9'b10000011;
				8'b1011110: c <= 9'b110000101;
				8'b1100111: c <= 9'b101101000;
				8'b1011010: c <= 9'b10101011;
				8'b1000010: c <= 9'b1010001;
				8'b111101: c <= 9'b100;
				8'b110000: c <= 9'b10110;
				8'b111110: c <= 9'b110100;
				8'b1100010: c <= 9'b100100000;
				8'b1110000: c <= 9'b111000111;
				8'b1101001: c <= 9'b101101001;
				8'b1110011: c <= 9'b110010111;
				8'b1001100: c <= 9'b100010101;
				8'b100001: c <= 9'b11101101;
				8'b1000110: c <= 9'b100010011;
				8'b1110010: c <= 9'b11111011;
				8'b1010000: c <= 9'b110110111;
				8'b1111010: c <= 9'b10100010;
				8'b1010101: c <= 9'b111110011;
				8'b111011: c <= 9'b100110101;
				8'b1001101: c <= 9'b100111;
				8'b111111: c <= 9'b1001101;
				8'b1101110: c <= 9'b10000010;
				8'b1111011: c <= 9'b1111010;
				8'b1001011: c <= 9'b1001101;
				8'b1101111: c <= 9'b110001010;
				8'b1101000: c <= 9'b101001001;
				8'b101100: c <= 9'b1000111;
				8'b100100: c <= 9'b1001100;
				8'b1111000: c <= 9'b110101100;
				8'b1000101: c <= 9'b111001011;
				8'b1011001: c <= 9'b110000110;
				8'b110100: c <= 9'b11111101;
				8'b1111001: c <= 9'b110011111;
				8'b1110001: c <= 9'b1011111;
				8'b1001111: c <= 9'b101111000;
				8'b1100101: c <= 9'b100011;
				8'b1111110: c <= 9'b100111110;
				8'b1111100: c <= 9'b11010101;
				8'b1010110: c <= 9'b11111011;
				8'b110010: c <= 9'b100100000;
				8'b1101101: c <= 9'b1000101;
				8'b100011: c <= 9'b1000010;
				8'b1110101: c <= 9'b1101101;
				8'b1111101: c <= 9'b111101111;
				8'b101001: c <= 9'b11;
				8'b1010010: c <= 9'b111000;
				8'b1011000: c <= 9'b11011110;
				8'b101110: c <= 9'b100111110;
				8'b1000001: c <= 9'b101010010;
				default: c <= 9'b0;
			endcase
			9'b10100 : case(di)
				8'b1000011: c <= 9'b111011001;
				8'b101000: c <= 9'b111000101;
				8'b111010: c <= 9'b101110010;
				8'b110110: c <= 9'b100001101;
				8'b1100100: c <= 9'b10010001;
				8'b1000000: c <= 9'b111011111;
				8'b1110110: c <= 9'b1001001;
				8'b100101: c <= 9'b100011;
				8'b101111: c <= 9'b110011111;
				8'b100110: c <= 9'b10011000;
				8'b1100011: c <= 9'b11000001;
				8'b1001000: c <= 9'b10011010;
				8'b111000: c <= 9'b1101100;
				8'b110001: c <= 9'b101101010;
				8'b1010111: c <= 9'b101000011;
				8'b1001110: c <= 9'b11000010;
				8'b1101010: c <= 9'b1000111;
				8'b1001001: c <= 9'b111010111;
				8'b1100000: c <= 9'b1011110;
				8'b110111: c <= 9'b110100000;
				8'b1011101: c <= 9'b101011001;
				8'b1011011: c <= 9'b10100011;
				8'b111001: c <= 9'b101101000;
				8'b1001010: c <= 9'b100010001;
				8'b110011: c <= 9'b111000110;
				8'b1101100: c <= 9'b10010000;
				8'b1110111: c <= 9'b100110110;
				8'b101011: c <= 9'b110110000;
				8'b1101011: c <= 9'b101001010;
				8'b111100: c <= 9'b10010111;
				8'b1000111: c <= 9'b100011101;
				8'b1011111: c <= 9'b1001101;
				8'b1110100: c <= 9'b101100000;
				8'b101101: c <= 9'b10001000;
				8'b1010011: c <= 9'b100000111;
				8'b1100001: c <= 9'b101001100;
				8'b110101: c <= 9'b10110;
				8'b1000100: c <= 9'b101011010;
				8'b1010001: c <= 9'b100100101;
				8'b1010100: c <= 9'b10010001;
				8'b1100110: c <= 9'b10011111;
				8'b101010: c <= 9'b110000001;
				8'b1011110: c <= 9'b1101111;
				8'b1100111: c <= 9'b100110010;
				8'b1011010: c <= 9'b100101110;
				8'b1000010: c <= 9'b110100000;
				8'b111101: c <= 9'b111011011;
				8'b110000: c <= 9'b11100000;
				8'b111110: c <= 9'b1001000;
				8'b1100010: c <= 9'b11001100;
				8'b1110000: c <= 9'b100100011;
				8'b1101001: c <= 9'b110101110;
				8'b1110011: c <= 9'b101111001;
				8'b1001100: c <= 9'b1011111;
				8'b100001: c <= 9'b101111110;
				8'b1000110: c <= 9'b111100110;
				8'b1110010: c <= 9'b11110010;
				8'b1010000: c <= 9'b10000101;
				8'b1111010: c <= 9'b11100010;
				8'b1010101: c <= 9'b100100010;
				8'b111011: c <= 9'b101110100;
				8'b1001101: c <= 9'b101000101;
				8'b111111: c <= 9'b100010100;
				8'b1101110: c <= 9'b100101001;
				8'b1111011: c <= 9'b100101011;
				8'b1001011: c <= 9'b100000011;
				8'b1101111: c <= 9'b110010;
				8'b1101000: c <= 9'b110100000;
				8'b101100: c <= 9'b101100;
				8'b100100: c <= 9'b11110100;
				8'b1111000: c <= 9'b100011001;
				8'b1000101: c <= 9'b101110101;
				8'b1011001: c <= 9'b110111110;
				8'b110100: c <= 9'b101000011;
				8'b1111001: c <= 9'b100100111;
				8'b1110001: c <= 9'b100010011;
				8'b1001111: c <= 9'b10110110;
				8'b1100101: c <= 9'b10010101;
				8'b1111110: c <= 9'b11101001;
				8'b1111100: c <= 9'b10010111;
				8'b1010110: c <= 9'b111010110;
				8'b110010: c <= 9'b110010011;
				8'b1101101: c <= 9'b101011011;
				8'b100011: c <= 9'b10010101;
				8'b1110101: c <= 9'b110111;
				8'b1111101: c <= 9'b1000111;
				8'b101001: c <= 9'b111010000;
				8'b1010010: c <= 9'b111101100;
				8'b1011000: c <= 9'b110000001;
				8'b101110: c <= 9'b101001010;
				8'b1000001: c <= 9'b10010011;
				default: c <= 9'b0;
			endcase
			9'b100110111 : case(di)
				8'b1000011: c <= 9'b11010010;
				8'b101000: c <= 9'b10000001;
				8'b111010: c <= 9'b101010011;
				8'b110110: c <= 9'b101101101;
				8'b1100100: c <= 9'b100110;
				8'b1000000: c <= 9'b110001101;
				8'b1110110: c <= 9'b111101000;
				8'b100101: c <= 9'b101000010;
				8'b101111: c <= 9'b1011110;
				8'b100110: c <= 9'b1110101;
				8'b1100011: c <= 9'b10011;
				8'b1001000: c <= 9'b110000;
				8'b111000: c <= 9'b100011000;
				8'b110001: c <= 9'b110010110;
				8'b1010111: c <= 9'b100101010;
				8'b1001110: c <= 9'b10001111;
				8'b1101010: c <= 9'b10011011;
				8'b1001001: c <= 9'b10111000;
				8'b1100000: c <= 9'b10001000;
				8'b110111: c <= 9'b111100011;
				8'b1011101: c <= 9'b100;
				8'b1011011: c <= 9'b100010010;
				8'b111001: c <= 9'b111111001;
				8'b1001010: c <= 9'b111100000;
				8'b110011: c <= 9'b1010110;
				8'b1101100: c <= 9'b101101000;
				8'b1110111: c <= 9'b111011100;
				8'b101011: c <= 9'b101100001;
				8'b1101011: c <= 9'b11011100;
				8'b111100: c <= 9'b111010000;
				8'b1000111: c <= 9'b111100000;
				8'b1011111: c <= 9'b110011000;
				8'b1110100: c <= 9'b10101000;
				8'b101101: c <= 9'b1010010;
				8'b1010011: c <= 9'b110100;
				8'b1100001: c <= 9'b111100100;
				8'b110101: c <= 9'b101101;
				8'b1000100: c <= 9'b11010;
				8'b1010001: c <= 9'b110110011;
				8'b1010100: c <= 9'b100011000;
				8'b1100110: c <= 9'b110001100;
				8'b101010: c <= 9'b110001;
				8'b1011110: c <= 9'b11000100;
				8'b1100111: c <= 9'b10000111;
				8'b1011010: c <= 9'b111100111;
				8'b1000010: c <= 9'b100010011;
				8'b111101: c <= 9'b101000001;
				8'b110000: c <= 9'b100010110;
				8'b111110: c <= 9'b100010000;
				8'b1100010: c <= 9'b1111;
				8'b1110000: c <= 9'b1001;
				8'b1101001: c <= 9'b111111000;
				8'b1110011: c <= 9'b111010;
				8'b1001100: c <= 9'b101011101;
				8'b100001: c <= 9'b10010110;
				8'b1000110: c <= 9'b111110011;
				8'b1110010: c <= 9'b100001101;
				8'b1010000: c <= 9'b100010010;
				8'b1111010: c <= 9'b101110100;
				8'b1010101: c <= 9'b100111000;
				8'b111011: c <= 9'b111000000;
				8'b1001101: c <= 9'b10111101;
				8'b111111: c <= 9'b100111010;
				8'b1101110: c <= 9'b111010111;
				8'b1111011: c <= 9'b101101001;
				8'b1001011: c <= 9'b110011010;
				8'b1101111: c <= 9'b101100100;
				8'b1101000: c <= 9'b111100;
				8'b101100: c <= 9'b100011;
				8'b100100: c <= 9'b100011001;
				8'b1111000: c <= 9'b101101110;
				8'b1000101: c <= 9'b11110;
				8'b1011001: c <= 9'b100010100;
				8'b110100: c <= 9'b10110111;
				8'b1111001: c <= 9'b110101;
				8'b1110001: c <= 9'b11110000;
				8'b1001111: c <= 9'b1101010;
				8'b1100101: c <= 9'b110101101;
				8'b1111110: c <= 9'b100001110;
				8'b1111100: c <= 9'b100011101;
				8'b1010110: c <= 9'b1101101;
				8'b110010: c <= 9'b111100;
				8'b1101101: c <= 9'b110000000;
				8'b100011: c <= 9'b110001;
				8'b1110101: c <= 9'b11000011;
				8'b1111101: c <= 9'b111110011;
				8'b101001: c <= 9'b10010111;
				8'b1010010: c <= 9'b110010001;
				8'b1011000: c <= 9'b1110011;
				8'b101110: c <= 9'b11000110;
				8'b1000001: c <= 9'b101111111;
				default: c <= 9'b0;
			endcase
			9'b110011100 : case(di)
				8'b1000011: c <= 9'b110010100;
				8'b101000: c <= 9'b11101011;
				8'b111010: c <= 9'b100111;
				8'b110110: c <= 9'b110101111;
				8'b1100100: c <= 9'b111000101;
				8'b1000000: c <= 9'b110111011;
				8'b1110110: c <= 9'b110011001;
				8'b100101: c <= 9'b110101111;
				8'b101111: c <= 9'b110010100;
				8'b100110: c <= 9'b100100111;
				8'b1100011: c <= 9'b1011001;
				8'b1001000: c <= 9'b100010011;
				8'b111000: c <= 9'b100100;
				8'b110001: c <= 9'b111010;
				8'b1010111: c <= 9'b10001010;
				8'b1001110: c <= 9'b11110110;
				8'b1101010: c <= 9'b111000;
				8'b1001001: c <= 9'b101111000;
				8'b1100000: c <= 9'b100000110;
				8'b110111: c <= 9'b11111;
				8'b1011101: c <= 9'b1010011;
				8'b1011011: c <= 9'b110101001;
				8'b111001: c <= 9'b100111010;
				8'b1001010: c <= 9'b1111001;
				8'b110011: c <= 9'b1101100;
				8'b1101100: c <= 9'b10001000;
				8'b1110111: c <= 9'b11;
				8'b101011: c <= 9'b110;
				8'b1101011: c <= 9'b11001000;
				8'b111100: c <= 9'b111011;
				8'b1000111: c <= 9'b1000111;
				8'b1011111: c <= 9'b1011011;
				8'b1110100: c <= 9'b110001000;
				8'b101101: c <= 9'b100110000;
				8'b1010011: c <= 9'b11000110;
				8'b1100001: c <= 9'b110000111;
				8'b110101: c <= 9'b11111010;
				8'b1000100: c <= 9'b111101111;
				8'b1010001: c <= 9'b10000000;
				8'b1010100: c <= 9'b111100010;
				8'b1100110: c <= 9'b100110111;
				8'b101010: c <= 9'b111110011;
				8'b1011110: c <= 9'b1000110;
				8'b1100111: c <= 9'b110010111;
				8'b1011010: c <= 9'b110011100;
				8'b1000010: c <= 9'b11110101;
				8'b111101: c <= 9'b1110100;
				8'b110000: c <= 9'b100111000;
				8'b111110: c <= 9'b110001111;
				8'b1100010: c <= 9'b110011001;
				8'b1110000: c <= 9'b101010000;
				8'b1101001: c <= 9'b1111;
				8'b1110011: c <= 9'b10000000;
				8'b1001100: c <= 9'b1010110;
				8'b100001: c <= 9'b10100;
				8'b1000110: c <= 9'b110001110;
				8'b1110010: c <= 9'b101010010;
				8'b1010000: c <= 9'b100011101;
				8'b1111010: c <= 9'b110011100;
				8'b1010101: c <= 9'b110111110;
				8'b111011: c <= 9'b10111001;
				8'b1001101: c <= 9'b101;
				8'b111111: c <= 9'b110010101;
				8'b1101110: c <= 9'b111001110;
				8'b1111011: c <= 9'b110000010;
				8'b1001011: c <= 9'b11001111;
				8'b1101111: c <= 9'b101010001;
				8'b1101000: c <= 9'b101010001;
				8'b101100: c <= 9'b111000101;
				8'b100100: c <= 9'b101110110;
				8'b1111000: c <= 9'b10101;
				8'b1000101: c <= 9'b100111001;
				8'b1011001: c <= 9'b110101010;
				8'b110100: c <= 9'b111100000;
				8'b1111001: c <= 9'b101110;
				8'b1110001: c <= 9'b1110111;
				8'b1001111: c <= 9'b110100;
				8'b1100101: c <= 9'b1001010;
				8'b1111110: c <= 9'b101101101;
				8'b1111100: c <= 9'b110001;
				8'b1010110: c <= 9'b10101;
				8'b110010: c <= 9'b111110101;
				8'b1101101: c <= 9'b100110101;
				8'b100011: c <= 9'b11010;
				8'b1110101: c <= 9'b111011010;
				8'b1111101: c <= 9'b111010111;
				8'b101001: c <= 9'b1111000;
				8'b1010010: c <= 9'b11010010;
				8'b1011000: c <= 9'b10000011;
				8'b101110: c <= 9'b110001111;
				8'b1000001: c <= 9'b10110011;
				default: c <= 9'b0;
			endcase
			9'b100001110 : case(di)
				8'b1000011: c <= 9'b100100101;
				8'b101000: c <= 9'b1110001;
				8'b111010: c <= 9'b11010100;
				8'b110110: c <= 9'b111010001;
				8'b1100100: c <= 9'b110010011;
				8'b1000000: c <= 9'b11000010;
				8'b1110110: c <= 9'b1100000;
				8'b100101: c <= 9'b11010101;
				8'b101111: c <= 9'b10000010;
				8'b100110: c <= 9'b10100000;
				8'b1100011: c <= 9'b10100110;
				8'b1001000: c <= 9'b11100100;
				8'b111000: c <= 9'b110011001;
				8'b110001: c <= 9'b1010001;
				8'b1010111: c <= 9'b1111110;
				8'b1001110: c <= 9'b1100011;
				8'b1101010: c <= 9'b1111110;
				8'b1001001: c <= 9'b11100101;
				8'b1100000: c <= 9'b111001111;
				8'b110111: c <= 9'b10000110;
				8'b1011101: c <= 9'b100111101;
				8'b1011011: c <= 9'b100011000;
				8'b111001: c <= 9'b110101010;
				8'b1001010: c <= 9'b110101001;
				8'b110011: c <= 9'b11101000;
				8'b1101100: c <= 9'b1100011;
				8'b1110111: c <= 9'b110010100;
				8'b101011: c <= 9'b101010;
				8'b1101011: c <= 9'b10101111;
				8'b111100: c <= 9'b100101;
				8'b1000111: c <= 9'b110100001;
				8'b1011111: c <= 9'b100111010;
				8'b1110100: c <= 9'b111011001;
				8'b101101: c <= 9'b1011001;
				8'b1010011: c <= 9'b100001;
				8'b1100001: c <= 9'b10001110;
				8'b110101: c <= 9'b10010;
				8'b1000100: c <= 9'b111000100;
				8'b1010001: c <= 9'b110111110;
				8'b1010100: c <= 9'b11111101;
				8'b1100110: c <= 9'b101011110;
				8'b101010: c <= 9'b101000001;
				8'b1011110: c <= 9'b101100100;
				8'b1100111: c <= 9'b111011001;
				8'b1011010: c <= 9'b110100100;
				8'b1000010: c <= 9'b100100011;
				8'b111101: c <= 9'b11000010;
				8'b110000: c <= 9'b101100000;
				8'b111110: c <= 9'b11111100;
				8'b1100010: c <= 9'b10000000;
				8'b1110000: c <= 9'b111000011;
				8'b1101001: c <= 9'b1010001;
				8'b1110011: c <= 9'b1000;
				8'b1001100: c <= 9'b110000010;
				8'b100001: c <= 9'b10000101;
				8'b1000110: c <= 9'b11111000;
				8'b1110010: c <= 9'b110111011;
				8'b1010000: c <= 9'b100000011;
				8'b1111010: c <= 9'b100001111;
				8'b1010101: c <= 9'b101100111;
				8'b111011: c <= 9'b11101011;
				8'b1001101: c <= 9'b111001;
				8'b111111: c <= 9'b10011000;
				8'b1101110: c <= 9'b11010011;
				8'b1111011: c <= 9'b100110100;
				8'b1001011: c <= 9'b100000001;
				8'b1101111: c <= 9'b111001010;
				8'b1101000: c <= 9'b101010101;
				8'b101100: c <= 9'b110111;
				8'b100100: c <= 9'b101111010;
				8'b1111000: c <= 9'b101001011;
				8'b1000101: c <= 9'b10100000;
				8'b1011001: c <= 9'b100111;
				8'b110100: c <= 9'b1111110;
				8'b1111001: c <= 9'b110111;
				8'b1110001: c <= 9'b11000100;
				8'b1001111: c <= 9'b1001101;
				8'b1100101: c <= 9'b110011001;
				8'b1111110: c <= 9'b101001;
				8'b1111100: c <= 9'b110101;
				8'b1010110: c <= 9'b10110010;
				8'b110010: c <= 9'b110000000;
				8'b1101101: c <= 9'b11001100;
				8'b100011: c <= 9'b100001111;
				8'b1110101: c <= 9'b110100011;
				8'b1111101: c <= 9'b10000001;
				8'b101001: c <= 9'b100011;
				8'b1010010: c <= 9'b10110111;
				8'b1011000: c <= 9'b111100101;
				8'b101110: c <= 9'b101101111;
				8'b1000001: c <= 9'b111111111;
				default: c <= 9'b0;
			endcase
			9'b1101110 : case(di)
				8'b1000011: c <= 9'b110100111;
				8'b101000: c <= 9'b100011111;
				8'b111010: c <= 9'b111000010;
				8'b110110: c <= 9'b101111010;
				8'b1100100: c <= 9'b1011;
				8'b1000000: c <= 9'b11111010;
				8'b1110110: c <= 9'b110100100;
				8'b100101: c <= 9'b1101111;
				8'b101111: c <= 9'b10111111;
				8'b100110: c <= 9'b1000110;
				8'b1100011: c <= 9'b1001;
				8'b1001000: c <= 9'b110011111;
				8'b111000: c <= 9'b1010011;
				8'b110001: c <= 9'b101010;
				8'b1010111: c <= 9'b100001110;
				8'b1001110: c <= 9'b10101010;
				8'b1101010: c <= 9'b11000;
				8'b1001001: c <= 9'b10001000;
				8'b1100000: c <= 9'b101101010;
				8'b110111: c <= 9'b101010101;
				8'b1011101: c <= 9'b10111110;
				8'b1011011: c <= 9'b101100;
				8'b111001: c <= 9'b100100111;
				8'b1001010: c <= 9'b11010101;
				8'b110011: c <= 9'b11010011;
				8'b1101100: c <= 9'b1111010;
				8'b1110111: c <= 9'b1110001;
				8'b101011: c <= 9'b111110001;
				8'b1101011: c <= 9'b111011110;
				8'b111100: c <= 9'b110001010;
				8'b1000111: c <= 9'b11001010;
				8'b1011111: c <= 9'b1011011;
				8'b1110100: c <= 9'b111100110;
				8'b101101: c <= 9'b11010;
				8'b1010011: c <= 9'b110000101;
				8'b1100001: c <= 9'b100010111;
				8'b110101: c <= 9'b111000111;
				8'b1000100: c <= 9'b10110111;
				8'b1010001: c <= 9'b111101001;
				8'b1010100: c <= 9'b111010110;
				8'b1100110: c <= 9'b111101010;
				8'b101010: c <= 9'b101111111;
				8'b1011110: c <= 9'b100011100;
				8'b1100111: c <= 9'b101001;
				8'b1011010: c <= 9'b1110001;
				8'b1000010: c <= 9'b1100100;
				8'b111101: c <= 9'b110110110;
				8'b110000: c <= 9'b11100100;
				8'b111110: c <= 9'b100100110;
				8'b1100010: c <= 9'b11111;
				8'b1110000: c <= 9'b100000101;
				8'b1101001: c <= 9'b111000000;
				8'b1110011: c <= 9'b111101101;
				8'b1001100: c <= 9'b1110010;
				8'b100001: c <= 9'b101101111;
				8'b1000110: c <= 9'b11001;
				8'b1110010: c <= 9'b110110111;
				8'b1010000: c <= 9'b111111110;
				8'b1111010: c <= 9'b110101001;
				8'b1010101: c <= 9'b110011;
				8'b111011: c <= 9'b101010100;
				8'b1001101: c <= 9'b10111110;
				8'b111111: c <= 9'b1110111;
				8'b1101110: c <= 9'b11100100;
				8'b1111011: c <= 9'b111011001;
				8'b1001011: c <= 9'b100001111;
				8'b1101111: c <= 9'b1000;
				8'b1101000: c <= 9'b110011000;
				8'b101100: c <= 9'b111;
				8'b100100: c <= 9'b11111;
				8'b1111000: c <= 9'b1100011;
				8'b1000101: c <= 9'b11100111;
				8'b1011001: c <= 9'b100011111;
				8'b110100: c <= 9'b11011100;
				8'b1111001: c <= 9'b110110110;
				8'b1110001: c <= 9'b11010100;
				8'b1001111: c <= 9'b101011110;
				8'b1100101: c <= 9'b111111000;
				8'b1111110: c <= 9'b110110101;
				8'b1111100: c <= 9'b10011100;
				8'b1010110: c <= 9'b1001010;
				8'b110010: c <= 9'b10010;
				8'b1101101: c <= 9'b1000100;
				8'b100011: c <= 9'b10111010;
				8'b1110101: c <= 9'b101011011;
				8'b1111101: c <= 9'b110110110;
				8'b101001: c <= 9'b101101110;
				8'b1010010: c <= 9'b101101100;
				8'b1011000: c <= 9'b101000010;
				8'b101110: c <= 9'b111100001;
				8'b1000001: c <= 9'b1010010;
				default: c <= 9'b0;
			endcase
			9'b101011010 : case(di)
				8'b1000011: c <= 9'b100001010;
				8'b101000: c <= 9'b10111100;
				8'b111010: c <= 9'b100011111;
				8'b110110: c <= 9'b101110100;
				8'b1100100: c <= 9'b111010110;
				8'b1000000: c <= 9'b101011110;
				8'b1110110: c <= 9'b100111110;
				8'b100101: c <= 9'b101000010;
				8'b101111: c <= 9'b100010000;
				8'b100110: c <= 9'b10100110;
				8'b1100011: c <= 9'b100100101;
				8'b1001000: c <= 9'b1001101;
				8'b111000: c <= 9'b1110111;
				8'b110001: c <= 9'b11101100;
				8'b1010111: c <= 9'b101110000;
				8'b1001110: c <= 9'b110110000;
				8'b1101010: c <= 9'b110011;
				8'b1001001: c <= 9'b1010101;
				8'b1100000: c <= 9'b10010;
				8'b110111: c <= 9'b100110111;
				8'b1011101: c <= 9'b11001000;
				8'b1011011: c <= 9'b110100100;
				8'b111001: c <= 9'b11111;
				8'b1001010: c <= 9'b101011010;
				8'b110011: c <= 9'b1011111;
				8'b1101100: c <= 9'b1100001;
				8'b1110111: c <= 9'b1001101;
				8'b101011: c <= 9'b10011111;
				8'b1101011: c <= 9'b100010110;
				8'b111100: c <= 9'b1111000;
				8'b1000111: c <= 9'b10000101;
				8'b1011111: c <= 9'b111001;
				8'b1110100: c <= 9'b111110001;
				8'b101101: c <= 9'b1100001;
				8'b1010011: c <= 9'b110011101;
				8'b1100001: c <= 9'b101100100;
				8'b110101: c <= 9'b101101100;
				8'b1000100: c <= 9'b100101100;
				8'b1010001: c <= 9'b10010001;
				8'b1010100: c <= 9'b111111111;
				8'b1100110: c <= 9'b100100101;
				8'b101010: c <= 9'b100111111;
				8'b1011110: c <= 9'b110000010;
				8'b1100111: c <= 9'b11011;
				8'b1011010: c <= 9'b110001100;
				8'b1000010: c <= 9'b1100100;
				8'b111101: c <= 9'b111111000;
				8'b110000: c <= 9'b101100000;
				8'b111110: c <= 9'b110010100;
				8'b1100010: c <= 9'b10101110;
				8'b1110000: c <= 9'b110001000;
				8'b1101001: c <= 9'b111101101;
				8'b1110011: c <= 9'b100000010;
				8'b1001100: c <= 9'b111010;
				8'b100001: c <= 9'b110;
				8'b1000110: c <= 9'b11111011;
				8'b1110010: c <= 9'b101001110;
				8'b1010000: c <= 9'b110011010;
				8'b1111010: c <= 9'b1001001;
				8'b1010101: c <= 9'b101110000;
				8'b111011: c <= 9'b10111111;
				8'b1001101: c <= 9'b101101001;
				8'b111111: c <= 9'b111011;
				8'b1101110: c <= 9'b11010;
				8'b1111011: c <= 9'b111101001;
				8'b1001011: c <= 9'b101011111;
				8'b1101111: c <= 9'b10010;
				8'b1101000: c <= 9'b1001110;
				8'b101100: c <= 9'b1011001;
				8'b100100: c <= 9'b101011000;
				8'b1111000: c <= 9'b11101101;
				8'b1000101: c <= 9'b111001010;
				8'b1011001: c <= 9'b11101001;
				8'b110100: c <= 9'b11000011;
				8'b1111001: c <= 9'b110010001;
				8'b1110001: c <= 9'b100000000;
				8'b1001111: c <= 9'b110100011;
				8'b1100101: c <= 9'b10011001;
				8'b1111110: c <= 9'b10;
				8'b1111100: c <= 9'b1101000;
				8'b1010110: c <= 9'b1010001;
				8'b110010: c <= 9'b11001010;
				8'b1101101: c <= 9'b11111001;
				8'b100011: c <= 9'b110100000;
				8'b1110101: c <= 9'b11000000;
				8'b1111101: c <= 9'b111111010;
				8'b101001: c <= 9'b10011001;
				8'b1010010: c <= 9'b100011010;
				8'b1011000: c <= 9'b11100000;
				8'b101110: c <= 9'b110100010;
				8'b1000001: c <= 9'b10000010;
				default: c <= 9'b0;
			endcase
			9'b11100100 : case(di)
				8'b1000011: c <= 9'b111001111;
				8'b101000: c <= 9'b110;
				8'b111010: c <= 9'b100101000;
				8'b110110: c <= 9'b11100001;
				8'b1100100: c <= 9'b111111010;
				8'b1000000: c <= 9'b111010110;
				8'b1110110: c <= 9'b11001111;
				8'b100101: c <= 9'b100000111;
				8'b101111: c <= 9'b111001011;
				8'b100110: c <= 9'b110100100;
				8'b1100011: c <= 9'b10110100;
				8'b1001000: c <= 9'b10000011;
				8'b111000: c <= 9'b111101101;
				8'b110001: c <= 9'b1010011;
				8'b1010111: c <= 9'b11100000;
				8'b1001110: c <= 9'b100000100;
				8'b1101010: c <= 9'b10010110;
				8'b1001001: c <= 9'b11010001;
				8'b1100000: c <= 9'b1110;
				8'b110111: c <= 9'b11110101;
				8'b1011101: c <= 9'b11001110;
				8'b1011011: c <= 9'b110100001;
				8'b111001: c <= 9'b10011010;
				8'b1001010: c <= 9'b111100111;
				8'b110011: c <= 9'b1100;
				8'b1101100: c <= 9'b11011011;
				8'b1110111: c <= 9'b10011001;
				8'b101011: c <= 9'b110011000;
				8'b1101011: c <= 9'b1101010;
				8'b111100: c <= 9'b101000;
				8'b1000111: c <= 9'b10011111;
				8'b1011111: c <= 9'b10110100;
				8'b1110100: c <= 9'b101010111;
				8'b101101: c <= 9'b101001100;
				8'b1010011: c <= 9'b111101101;
				8'b1100001: c <= 9'b100100000;
				8'b110101: c <= 9'b10001010;
				8'b1000100: c <= 9'b110110101;
				8'b1010001: c <= 9'b1011110;
				8'b1010100: c <= 9'b101101000;
				8'b1100110: c <= 9'b110000111;
				8'b101010: c <= 9'b110100101;
				8'b1011110: c <= 9'b101110000;
				8'b1100111: c <= 9'b1100000;
				8'b1011010: c <= 9'b10111110;
				8'b1000010: c <= 9'b10000101;
				8'b111101: c <= 9'b111101010;
				8'b110000: c <= 9'b11000010;
				8'b111110: c <= 9'b100011111;
				8'b1100010: c <= 9'b111001011;
				8'b1110000: c <= 9'b100100110;
				8'b1101001: c <= 9'b110111010;
				8'b1110011: c <= 9'b100111100;
				8'b1001100: c <= 9'b1000;
				8'b100001: c <= 9'b101100111;
				8'b1000110: c <= 9'b111010000;
				8'b1110010: c <= 9'b10101011;
				8'b1010000: c <= 9'b100101101;
				8'b1111010: c <= 9'b101010011;
				8'b1010101: c <= 9'b1100001;
				8'b111011: c <= 9'b10101;
				8'b1001101: c <= 9'b10110;
				8'b111111: c <= 9'b111011110;
				8'b1101110: c <= 9'b1001101;
				8'b1111011: c <= 9'b100110111;
				8'b1001011: c <= 9'b11010111;
				8'b1101111: c <= 9'b110101;
				8'b1101000: c <= 9'b1101001;
				8'b101100: c <= 9'b100110;
				8'b100100: c <= 9'b100011111;
				8'b1111000: c <= 9'b10000010;
				8'b1000101: c <= 9'b11011100;
				8'b1011001: c <= 9'b101001010;
				8'b110100: c <= 9'b1010110;
				8'b1111001: c <= 9'b100111100;
				8'b1110001: c <= 9'b1001000;
				8'b1001111: c <= 9'b101101011;
				8'b1100101: c <= 9'b10101010;
				8'b1111110: c <= 9'b11100;
				8'b1111100: c <= 9'b1110011;
				8'b1010110: c <= 9'b100111001;
				8'b110010: c <= 9'b100100;
				8'b1101101: c <= 9'b100010000;
				8'b100011: c <= 9'b101110100;
				8'b1110101: c <= 9'b110000101;
				8'b1111101: c <= 9'b100001111;
				8'b101001: c <= 9'b110000010;
				8'b1010010: c <= 9'b111000010;
				8'b1011000: c <= 9'b100101110;
				8'b101110: c <= 9'b100110;
				8'b1000001: c <= 9'b100000001;
				default: c <= 9'b0;
			endcase
			9'b111001100 : case(di)
				8'b1000011: c <= 9'b111001101;
				8'b101000: c <= 9'b110001001;
				8'b111010: c <= 9'b110101001;
				8'b110110: c <= 9'b1101110;
				8'b1100100: c <= 9'b1111100;
				8'b1000000: c <= 9'b1010110;
				8'b1110110: c <= 9'b110010001;
				8'b100101: c <= 9'b110011001;
				8'b101111: c <= 9'b101001;
				8'b100110: c <= 9'b10000;
				8'b1100011: c <= 9'b110101110;
				8'b1001000: c <= 9'b100111010;
				8'b111000: c <= 9'b110100001;
				8'b110001: c <= 9'b110011;
				8'b1010111: c <= 9'b110001111;
				8'b1001110: c <= 9'b1011001;
				8'b1101010: c <= 9'b110001100;
				8'b1001001: c <= 9'b101001000;
				8'b1100000: c <= 9'b100110011;
				8'b110111: c <= 9'b101101110;
				8'b1011101: c <= 9'b1001101;
				8'b1011011: c <= 9'b100011011;
				8'b111001: c <= 9'b110101010;
				8'b1001010: c <= 9'b1010010;
				8'b110011: c <= 9'b110100;
				8'b1101100: c <= 9'b10111100;
				8'b1110111: c <= 9'b100001010;
				8'b101011: c <= 9'b1010000;
				8'b1101011: c <= 9'b10011010;
				8'b111100: c <= 9'b100101000;
				8'b1000111: c <= 9'b101000110;
				8'b1011111: c <= 9'b111011101;
				8'b1110100: c <= 9'b111110000;
				8'b101101: c <= 9'b111000011;
				8'b1010011: c <= 9'b111010;
				8'b1100001: c <= 9'b11000000;
				8'b110101: c <= 9'b110001001;
				8'b1000100: c <= 9'b110001001;
				8'b1010001: c <= 9'b110111;
				8'b1010100: c <= 9'b111101010;
				8'b1100110: c <= 9'b110010;
				8'b101010: c <= 9'b110100101;
				8'b1011110: c <= 9'b111101000;
				8'b1100111: c <= 9'b110110011;
				8'b1011010: c <= 9'b101001010;
				8'b1000010: c <= 9'b11110001;
				8'b111101: c <= 9'b11000111;
				8'b110000: c <= 9'b1101010;
				8'b111110: c <= 9'b11101111;
				8'b1100010: c <= 9'b101111110;
				8'b1110000: c <= 9'b111011100;
				8'b1101001: c <= 9'b100011010;
				8'b1110011: c <= 9'b111011110;
				8'b1001100: c <= 9'b110100011;
				8'b100001: c <= 9'b1111111;
				8'b1000110: c <= 9'b101010000;
				8'b1110010: c <= 9'b101110100;
				8'b1010000: c <= 9'b10100010;
				8'b1111010: c <= 9'b111000010;
				8'b1010101: c <= 9'b11100001;
				8'b111011: c <= 9'b110011101;
				8'b1001101: c <= 9'b11100111;
				8'b111111: c <= 9'b100010010;
				8'b1101110: c <= 9'b101011110;
				8'b1111011: c <= 9'b1100;
				8'b1001011: c <= 9'b100010010;
				8'b1101111: c <= 9'b11111010;
				8'b1101000: c <= 9'b111010000;
				8'b101100: c <= 9'b100001100;
				8'b100100: c <= 9'b1001110;
				8'b1111000: c <= 9'b1011010;
				8'b1000101: c <= 9'b1111011;
				8'b1011001: c <= 9'b110110101;
				8'b110100: c <= 9'b11000000;
				8'b1111001: c <= 9'b101011011;
				8'b1110001: c <= 9'b111110110;
				8'b1001111: c <= 9'b101010011;
				8'b1100101: c <= 9'b110010010;
				8'b1111110: c <= 9'b111111000;
				8'b1111100: c <= 9'b11010;
				8'b1010110: c <= 9'b10011010;
				8'b110010: c <= 9'b111011001;
				8'b1101101: c <= 9'b100010100;
				8'b100011: c <= 9'b101001000;
				8'b1110101: c <= 9'b1110000;
				8'b1111101: c <= 9'b111001101;
				8'b101001: c <= 9'b10110110;
				8'b1010010: c <= 9'b110110000;
				8'b1011000: c <= 9'b100101010;
				8'b101110: c <= 9'b1011;
				8'b1000001: c <= 9'b110010010;
				default: c <= 9'b0;
			endcase
			9'b10110110 : case(di)
				8'b1000011: c <= 9'b10010000;
				8'b101000: c <= 9'b10011010;
				8'b111010: c <= 9'b11011000;
				8'b110110: c <= 9'b1101100;
				8'b1100100: c <= 9'b100000101;
				8'b1000000: c <= 9'b11110000;
				8'b1110110: c <= 9'b101100100;
				8'b100101: c <= 9'b1001100;
				8'b101111: c <= 9'b10000111;
				8'b100110: c <= 9'b110011011;
				8'b1100011: c <= 9'b101010011;
				8'b1001000: c <= 9'b100110010;
				8'b111000: c <= 9'b11000;
				8'b110001: c <= 9'b101010000;
				8'b1010111: c <= 9'b111000111;
				8'b1001110: c <= 9'b111101000;
				8'b1101010: c <= 9'b11101;
				8'b1001001: c <= 9'b100011001;
				8'b1100000: c <= 9'b111001;
				8'b110111: c <= 9'b110011;
				8'b1011101: c <= 9'b110011011;
				8'b1011011: c <= 9'b1001010;
				8'b111001: c <= 9'b10000101;
				8'b1001010: c <= 9'b110000111;
				8'b110011: c <= 9'b101011110;
				8'b1101100: c <= 9'b1101100;
				8'b1110111: c <= 9'b1011010;
				8'b101011: c <= 9'b110010101;
				8'b1101011: c <= 9'b111;
				8'b111100: c <= 9'b111001;
				8'b1000111: c <= 9'b110011010;
				8'b1011111: c <= 9'b111000000;
				8'b1110100: c <= 9'b11010000;
				8'b101101: c <= 9'b100100110;
				8'b1010011: c <= 9'b101110111;
				8'b1100001: c <= 9'b1000011;
				8'b110101: c <= 9'b110010010;
				8'b1000100: c <= 9'b111101001;
				8'b1010001: c <= 9'b111001100;
				8'b1010100: c <= 9'b110011110;
				8'b1100110: c <= 9'b110000111;
				8'b101010: c <= 9'b11100000;
				8'b1011110: c <= 9'b11001;
				8'b1100111: c <= 9'b100011;
				8'b1011010: c <= 9'b1101000;
				8'b1000010: c <= 9'b110101001;
				8'b111101: c <= 9'b10100000;
				8'b110000: c <= 9'b111011110;
				8'b111110: c <= 9'b110000111;
				8'b1100010: c <= 9'b1110101;
				8'b1110000: c <= 9'b1001000;
				8'b1101001: c <= 9'b110111000;
				8'b1110011: c <= 9'b110101;
				8'b1001100: c <= 9'b110101010;
				8'b100001: c <= 9'b11110000;
				8'b1000110: c <= 9'b10100100;
				8'b1110010: c <= 9'b101011;
				8'b1010000: c <= 9'b1000001;
				8'b1111010: c <= 9'b110001010;
				8'b1010101: c <= 9'b101;
				8'b111011: c <= 9'b1100011;
				8'b1001101: c <= 9'b11000110;
				8'b111111: c <= 9'b1101010;
				8'b1101110: c <= 9'b111111101;
				8'b1111011: c <= 9'b1000011;
				8'b1001011: c <= 9'b1101;
				8'b1101111: c <= 9'b100110;
				8'b1101000: c <= 9'b10111111;
				8'b101100: c <= 9'b100100111;
				8'b100100: c <= 9'b1101010;
				8'b1111000: c <= 9'b10100;
				8'b1000101: c <= 9'b110110101;
				8'b1011001: c <= 9'b11100101;
				8'b110100: c <= 9'b1010001;
				8'b1111001: c <= 9'b111011010;
				8'b1110001: c <= 9'b1000011;
				8'b1001111: c <= 9'b1100111;
				8'b1100101: c <= 9'b101;
				8'b1111110: c <= 9'b10001110;
				8'b1111100: c <= 9'b111110000;
				8'b1010110: c <= 9'b101101101;
				8'b110010: c <= 9'b100011010;
				8'b1101101: c <= 9'b11011010;
				8'b100011: c <= 9'b10100000;
				8'b1110101: c <= 9'b110010;
				8'b1111101: c <= 9'b1101110;
				8'b101001: c <= 9'b100110101;
				8'b1010010: c <= 9'b100000001;
				8'b1011000: c <= 9'b100001101;
				8'b101110: c <= 9'b11111010;
				8'b1000001: c <= 9'b100111100;
				default: c <= 9'b0;
			endcase
			9'b111101000 : case(di)
				8'b1000011: c <= 9'b111001101;
				8'b101000: c <= 9'b101101101;
				8'b111010: c <= 9'b1010001;
				8'b110110: c <= 9'b100101001;
				8'b1100100: c <= 9'b101000011;
				8'b1000000: c <= 9'b1101010;
				8'b1110110: c <= 9'b11010101;
				8'b100101: c <= 9'b111100111;
				8'b101111: c <= 9'b100111101;
				8'b100110: c <= 9'b11000110;
				8'b1100011: c <= 9'b10001100;
				8'b1001000: c <= 9'b100011111;
				8'b111000: c <= 9'b10011111;
				8'b110001: c <= 9'b111001110;
				8'b1010111: c <= 9'b11000100;
				8'b1001110: c <= 9'b110111;
				8'b1101010: c <= 9'b11100001;
				8'b1001001: c <= 9'b101000;
				8'b1100000: c <= 9'b10011000;
				8'b110111: c <= 9'b1101000;
				8'b1011101: c <= 9'b111100001;
				8'b1011011: c <= 9'b11110010;
				8'b111001: c <= 9'b111101110;
				8'b1001010: c <= 9'b101001000;
				8'b110011: c <= 9'b1000011;
				8'b1101100: c <= 9'b11000010;
				8'b1110111: c <= 9'b110011100;
				8'b101011: c <= 9'b1010000;
				8'b1101011: c <= 9'b1;
				8'b111100: c <= 9'b11011101;
				8'b1000111: c <= 9'b100011;
				8'b1011111: c <= 9'b110111011;
				8'b1110100: c <= 9'b101110100;
				8'b101101: c <= 9'b111110001;
				8'b1010011: c <= 9'b101000101;
				8'b1100001: c <= 9'b111100110;
				8'b110101: c <= 9'b110111110;
				8'b1000100: c <= 9'b111111011;
				8'b1010001: c <= 9'b1000100;
				8'b1010100: c <= 9'b11011001;
				8'b1100110: c <= 9'b100011000;
				8'b101010: c <= 9'b100000101;
				8'b1011110: c <= 9'b11010000;
				8'b1100111: c <= 9'b111001101;
				8'b1011010: c <= 9'b111101;
				8'b1000010: c <= 9'b101010100;
				8'b111101: c <= 9'b110101;
				8'b110000: c <= 9'b10000010;
				8'b111110: c <= 9'b1011111;
				8'b1100010: c <= 9'b10111110;
				8'b1110000: c <= 9'b11100110;
				8'b1101001: c <= 9'b110110010;
				8'b1110011: c <= 9'b11011011;
				8'b1001100: c <= 9'b11110001;
				8'b100001: c <= 9'b10010100;
				8'b1000110: c <= 9'b10111;
				8'b1110010: c <= 9'b11010100;
				8'b1010000: c <= 9'b100111000;
				8'b1111010: c <= 9'b1100110;
				8'b1010101: c <= 9'b11010100;
				8'b111011: c <= 9'b1100100;
				8'b1001101: c <= 9'b111110110;
				8'b111111: c <= 9'b1101111;
				8'b1101110: c <= 9'b10010;
				8'b1111011: c <= 9'b110111111;
				8'b1001011: c <= 9'b111000010;
				8'b1101111: c <= 9'b11011110;
				8'b1101000: c <= 9'b111001101;
				8'b101100: c <= 9'b111010010;
				8'b100100: c <= 9'b1001110;
				8'b1111000: c <= 9'b11011;
				8'b1000101: c <= 9'b1010111;
				8'b1011001: c <= 9'b10001010;
				8'b110100: c <= 9'b110011101;
				8'b1111001: c <= 9'b1100011;
				8'b1110001: c <= 9'b110000;
				8'b1001111: c <= 9'b100011001;
				8'b1100101: c <= 9'b111110000;
				8'b1111110: c <= 9'b11001100;
				8'b1111100: c <= 9'b10010100;
				8'b1010110: c <= 9'b100000000;
				8'b110010: c <= 9'b100001010;
				8'b1101101: c <= 9'b110111010;
				8'b100011: c <= 9'b1001000;
				8'b1110101: c <= 9'b101011010;
				8'b1111101: c <= 9'b10111100;
				8'b101001: c <= 9'b111101;
				8'b1010010: c <= 9'b110000111;
				8'b1011000: c <= 9'b100001;
				8'b101110: c <= 9'b101101001;
				8'b1000001: c <= 9'b110111010;
				default: c <= 9'b0;
			endcase
			9'b1110101 : case(di)
				8'b1000011: c <= 9'b101100110;
				8'b101000: c <= 9'b111000010;
				8'b111010: c <= 9'b111110000;
				8'b110110: c <= 9'b101100010;
				8'b1100100: c <= 9'b100010;
				8'b1000000: c <= 9'b111101111;
				8'b1110110: c <= 9'b10111010;
				8'b100101: c <= 9'b11100110;
				8'b101111: c <= 9'b100010010;
				8'b100110: c <= 9'b1101000;
				8'b1100011: c <= 9'b1111000;
				8'b1001000: c <= 9'b1111111;
				8'b111000: c <= 9'b1000111;
				8'b110001: c <= 9'b10100;
				8'b1010111: c <= 9'b101111010;
				8'b1001110: c <= 9'b111001000;
				8'b1101010: c <= 9'b100011001;
				8'b1001001: c <= 9'b110100000;
				8'b1100000: c <= 9'b1010111;
				8'b110111: c <= 9'b10011010;
				8'b1011101: c <= 9'b101001001;
				8'b1011011: c <= 9'b1111010;
				8'b111001: c <= 9'b1111100;
				8'b1001010: c <= 9'b110111;
				8'b110011: c <= 9'b101011;
				8'b1101100: c <= 9'b10001000;
				8'b1110111: c <= 9'b10001111;
				8'b101011: c <= 9'b1011;
				8'b1101011: c <= 9'b110100011;
				8'b111100: c <= 9'b111100001;
				8'b1000111: c <= 9'b1001;
				8'b1011111: c <= 9'b111010;
				8'b1110100: c <= 9'b101101001;
				8'b101101: c <= 9'b101011000;
				8'b1010011: c <= 9'b11100110;
				8'b1100001: c <= 9'b101110111;
				8'b110101: c <= 9'b101000011;
				8'b1000100: c <= 9'b110100100;
				8'b1010001: c <= 9'b100001110;
				8'b1010100: c <= 9'b111000000;
				8'b1100110: c <= 9'b10101101;
				8'b101010: c <= 9'b1111;
				8'b1011110: c <= 9'b110100000;
				8'b1100111: c <= 9'b1001;
				8'b1011010: c <= 9'b100101011;
				8'b1000010: c <= 9'b110000101;
				8'b111101: c <= 9'b110010100;
				8'b110000: c <= 9'b11111110;
				8'b111110: c <= 9'b1100000;
				8'b1100010: c <= 9'b110101111;
				8'b1110000: c <= 9'b110001100;
				8'b1101001: c <= 9'b11001101;
				8'b1110011: c <= 9'b11100101;
				8'b1001100: c <= 9'b10001000;
				8'b100001: c <= 9'b100110101;
				8'b1000110: c <= 9'b101001001;
				8'b1110010: c <= 9'b1111111;
				8'b1010000: c <= 9'b111000110;
				8'b1111010: c <= 9'b11111101;
				8'b1010101: c <= 9'b111010000;
				8'b111011: c <= 9'b110100001;
				8'b1001101: c <= 9'b101111000;
				8'b111111: c <= 9'b100011101;
				8'b1101110: c <= 9'b111101000;
				8'b1111011: c <= 9'b111011110;
				8'b1001011: c <= 9'b100;
				8'b1101111: c <= 9'b1101100;
				8'b1101000: c <= 9'b110001011;
				8'b101100: c <= 9'b10101;
				8'b100100: c <= 9'b110000011;
				8'b1111000: c <= 9'b100010100;
				8'b1000101: c <= 9'b111010000;
				8'b1011001: c <= 9'b1001101;
				8'b110100: c <= 9'b10011011;
				8'b1111001: c <= 9'b10110101;
				8'b1110001: c <= 9'b101111000;
				8'b1001111: c <= 9'b101011111;
				8'b1100101: c <= 9'b11100011;
				8'b1111110: c <= 9'b100100010;
				8'b1111100: c <= 9'b11110111;
				8'b1010110: c <= 9'b10000001;
				8'b110010: c <= 9'b100111110;
				8'b1101101: c <= 9'b100011100;
				8'b100011: c <= 9'b1000110;
				8'b1110101: c <= 9'b1011000;
				8'b1111101: c <= 9'b1011010;
				8'b101001: c <= 9'b1111;
				8'b1010010: c <= 9'b11011110;
				8'b1011000: c <= 9'b100010100;
				8'b101110: c <= 9'b111011011;
				8'b1000001: c <= 9'b111100001;
				default: c <= 9'b0;
			endcase
			9'b111011011 : case(di)
				8'b1000011: c <= 9'b1111001;
				8'b101000: c <= 9'b10101000;
				8'b111010: c <= 9'b10100110;
				8'b110110: c <= 9'b111011111;
				8'b1100100: c <= 9'b110100011;
				8'b1000000: c <= 9'b101111110;
				8'b1110110: c <= 9'b11100110;
				8'b100101: c <= 9'b11110010;
				8'b101111: c <= 9'b100010000;
				8'b100110: c <= 9'b110101001;
				8'b1100011: c <= 9'b10100000;
				8'b1001000: c <= 9'b111010001;
				8'b111000: c <= 9'b11110010;
				8'b110001: c <= 9'b101111001;
				8'b1010111: c <= 9'b1110011;
				8'b1001110: c <= 9'b10110;
				8'b1101010: c <= 9'b10101010;
				8'b1001001: c <= 9'b10010100;
				8'b1100000: c <= 9'b100100101;
				8'b110111: c <= 9'b11011000;
				8'b1011101: c <= 9'b100011;
				8'b1011011: c <= 9'b110000110;
				8'b111001: c <= 9'b110010010;
				8'b1001010: c <= 9'b110001101;
				8'b110011: c <= 9'b100000010;
				8'b1101100: c <= 9'b101001111;
				8'b1110111: c <= 9'b11;
				8'b101011: c <= 9'b101010000;
				8'b1101011: c <= 9'b10110110;
				8'b111100: c <= 9'b1001010;
				8'b1000111: c <= 9'b111001;
				8'b1011111: c <= 9'b10110011;
				8'b1110100: c <= 9'b111000;
				8'b101101: c <= 9'b111010010;
				8'b1010011: c <= 9'b10001010;
				8'b1100001: c <= 9'b1100111;
				8'b110101: c <= 9'b10101011;
				8'b1000100: c <= 9'b111100111;
				8'b1010001: c <= 9'b100010010;
				8'b1010100: c <= 9'b111111110;
				8'b1100110: c <= 9'b100001001;
				8'b101010: c <= 9'b11111001;
				8'b1011110: c <= 9'b101110010;
				8'b1100111: c <= 9'b10110010;
				8'b1011010: c <= 9'b111100011;
				8'b1000010: c <= 9'b100000010;
				8'b111101: c <= 9'b10010001;
				8'b110000: c <= 9'b111001010;
				8'b111110: c <= 9'b101100010;
				8'b1100010: c <= 9'b101000101;
				8'b1110000: c <= 9'b111000101;
				8'b1101001: c <= 9'b10010111;
				8'b1110011: c <= 9'b101011111;
				8'b1001100: c <= 9'b1100000;
				8'b100001: c <= 9'b10111111;
				8'b1000110: c <= 9'b110110101;
				8'b1110010: c <= 9'b110110;
				8'b1010000: c <= 9'b100110100;
				8'b1111010: c <= 9'b110100000;
				8'b1010101: c <= 9'b110110;
				8'b111011: c <= 9'b100110000;
				8'b1001101: c <= 9'b11001001;
				8'b111111: c <= 9'b101100001;
				8'b1101110: c <= 9'b101110100;
				8'b1111011: c <= 9'b110001100;
				8'b1001011: c <= 9'b10000111;
				8'b1101111: c <= 9'b100010;
				8'b1101000: c <= 9'b11110000;
				8'b101100: c <= 9'b111100001;
				8'b100100: c <= 9'b110111;
				8'b1111000: c <= 9'b1001110;
				8'b1000101: c <= 9'b11001011;
				8'b1011001: c <= 9'b10111011;
				8'b110100: c <= 9'b100001011;
				8'b1111001: c <= 9'b110101110;
				8'b1110001: c <= 9'b10110;
				8'b1001111: c <= 9'b100111111;
				8'b1100101: c <= 9'b111000101;
				8'b1111110: c <= 9'b10100011;
				8'b1111100: c <= 9'b10011011;
				8'b1010110: c <= 9'b10010110;
				8'b110010: c <= 9'b101111111;
				8'b1101101: c <= 9'b1;
				8'b100011: c <= 9'b1011100;
				8'b1110101: c <= 9'b101010101;
				8'b1111101: c <= 9'b10000000;
				8'b101001: c <= 9'b10100011;
				8'b1010010: c <= 9'b10000110;
				8'b1011000: c <= 9'b10111101;
				8'b101110: c <= 9'b101000101;
				8'b1000001: c <= 9'b1100100;
				default: c <= 9'b0;
			endcase
			9'b110111010 : case(di)
				8'b1000011: c <= 9'b1010001;
				8'b101000: c <= 9'b10110;
				8'b111010: c <= 9'b10011;
				8'b110110: c <= 9'b11001;
				8'b1100100: c <= 9'b100111100;
				8'b1000000: c <= 9'b11111;
				8'b1110110: c <= 9'b111010000;
				8'b100101: c <= 9'b110010100;
				8'b101111: c <= 9'b1101101;
				8'b100110: c <= 9'b11011000;
				8'b1100011: c <= 9'b100110;
				8'b1001000: c <= 9'b110101001;
				8'b111000: c <= 9'b10111001;
				8'b110001: c <= 9'b11110010;
				8'b1010111: c <= 9'b11101100;
				8'b1001110: c <= 9'b11010100;
				8'b1101010: c <= 9'b101000111;
				8'b1001001: c <= 9'b110010100;
				8'b1100000: c <= 9'b111010110;
				8'b110111: c <= 9'b100011100;
				8'b1011101: c <= 9'b11000100;
				8'b1011011: c <= 9'b1111001;
				8'b111001: c <= 9'b10111011;
				8'b1001010: c <= 9'b110001100;
				8'b110011: c <= 9'b101001100;
				8'b1101100: c <= 9'b111010001;
				8'b1110111: c <= 9'b1011000;
				8'b101011: c <= 9'b11110011;
				8'b1101011: c <= 9'b100001001;
				8'b111100: c <= 9'b110000;
				8'b1000111: c <= 9'b1011000;
				8'b1011111: c <= 9'b101010011;
				8'b1110100: c <= 9'b1011011;
				8'b101101: c <= 9'b110011111;
				8'b1010011: c <= 9'b111111010;
				8'b1100001: c <= 9'b1101001;
				8'b110101: c <= 9'b10111110;
				8'b1000100: c <= 9'b10010011;
				8'b1010001: c <= 9'b111001111;
				8'b1010100: c <= 9'b110110101;
				8'b1100110: c <= 9'b1001101;
				8'b101010: c <= 9'b10101011;
				8'b1011110: c <= 9'b111001;
				8'b1100111: c <= 9'b1101001;
				8'b1011010: c <= 9'b111110001;
				8'b1000010: c <= 9'b11001010;
				8'b111101: c <= 9'b11111100;
				8'b110000: c <= 9'b110000000;
				8'b111110: c <= 9'b111000111;
				8'b1100010: c <= 9'b111010010;
				8'b1110000: c <= 9'b110101110;
				8'b1101001: c <= 9'b111111101;
				8'b1110011: c <= 9'b110000110;
				8'b1001100: c <= 9'b111011;
				8'b100001: c <= 9'b11001;
				8'b1000110: c <= 9'b100110100;
				8'b1110010: c <= 9'b1101;
				8'b1010000: c <= 9'b10011111;
				8'b1111010: c <= 9'b101100001;
				8'b1010101: c <= 9'b111000;
				8'b111011: c <= 9'b110010;
				8'b1001101: c <= 9'b101100000;
				8'b111111: c <= 9'b101111111;
				8'b1101110: c <= 9'b11010010;
				8'b1111011: c <= 9'b11010100;
				8'b1001011: c <= 9'b1001100;
				8'b1101111: c <= 9'b11100011;
				8'b1101000: c <= 9'b110111110;
				8'b101100: c <= 9'b1001111;
				8'b100100: c <= 9'b1101110;
				8'b1111000: c <= 9'b111010111;
				8'b1000101: c <= 9'b1001100;
				8'b1011001: c <= 9'b100110011;
				8'b110100: c <= 9'b101101111;
				8'b1111001: c <= 9'b11001101;
				8'b1110001: c <= 9'b11101011;
				8'b1001111: c <= 9'b10111000;
				8'b1100101: c <= 9'b101001110;
				8'b1111110: c <= 9'b110110;
				8'b1111100: c <= 9'b10110010;
				8'b1010110: c <= 9'b100001111;
				8'b110010: c <= 9'b110010010;
				8'b1101101: c <= 9'b11010010;
				8'b100011: c <= 9'b110111001;
				8'b1110101: c <= 9'b11110010;
				8'b1111101: c <= 9'b110101111;
				8'b101001: c <= 9'b100111000;
				8'b1010010: c <= 9'b111001110;
				8'b1011000: c <= 9'b101001001;
				8'b101110: c <= 9'b110100011;
				8'b1000001: c <= 9'b1110111;
				default: c <= 9'b0;
			endcase
			9'b111101001 : case(di)
				8'b1000011: c <= 9'b11001111;
				8'b101000: c <= 9'b100011;
				8'b111010: c <= 9'b100010001;
				8'b110110: c <= 9'b110101101;
				8'b1100100: c <= 9'b110101001;
				8'b1000000: c <= 9'b10100011;
				8'b1110110: c <= 9'b10100010;
				8'b100101: c <= 9'b101011010;
				8'b101111: c <= 9'b101011110;
				8'b100110: c <= 9'b11000;
				8'b1100011: c <= 9'b111010;
				8'b1001000: c <= 9'b11000110;
				8'b111000: c <= 9'b110000111;
				8'b110001: c <= 9'b11001111;
				8'b1010111: c <= 9'b100011000;
				8'b1001110: c <= 9'b10001010;
				8'b1101010: c <= 9'b11011101;
				8'b1001001: c <= 9'b110010011;
				8'b1100000: c <= 9'b10110101;
				8'b110111: c <= 9'b110011100;
				8'b1011101: c <= 9'b11001;
				8'b1011011: c <= 9'b110100;
				8'b111001: c <= 9'b1100;
				8'b1001010: c <= 9'b110001001;
				8'b110011: c <= 9'b1;
				8'b1101100: c <= 9'b1001111;
				8'b1110111: c <= 9'b1100101;
				8'b101011: c <= 9'b100000100;
				8'b1101011: c <= 9'b10100;
				8'b111100: c <= 9'b1010001;
				8'b1000111: c <= 9'b1111111;
				8'b1011111: c <= 9'b111111;
				8'b1110100: c <= 9'b10111111;
				8'b101101: c <= 9'b10101000;
				8'b1010011: c <= 9'b110101001;
				8'b1100001: c <= 9'b101111110;
				8'b110101: c <= 9'b11110011;
				8'b1000100: c <= 9'b10101001;
				8'b1010001: c <= 9'b100111000;
				8'b1010100: c <= 9'b111001011;
				8'b1100110: c <= 9'b100011100;
				8'b101010: c <= 9'b1011110;
				8'b1011110: c <= 9'b11110100;
				8'b1100111: c <= 9'b10101001;
				8'b1011010: c <= 9'b111100010;
				8'b1000010: c <= 9'b10001111;
				8'b111101: c <= 9'b101010110;
				8'b110000: c <= 9'b1001010;
				8'b111110: c <= 9'b110101;
				8'b1100010: c <= 9'b1000110;
				8'b1110000: c <= 9'b111011001;
				8'b1101001: c <= 9'b111011110;
				8'b1110011: c <= 9'b11101101;
				8'b1001100: c <= 9'b111011100;
				8'b100001: c <= 9'b101000111;
				8'b1000110: c <= 9'b11101111;
				8'b1110010: c <= 9'b1000100;
				8'b1010000: c <= 9'b10101001;
				8'b1111010: c <= 9'b1001000;
				8'b1010101: c <= 9'b110010010;
				8'b111011: c <= 9'b110000010;
				8'b1001101: c <= 9'b100100010;
				8'b111111: c <= 9'b10100010;
				8'b1101110: c <= 9'b10011010;
				8'b1111011: c <= 9'b11010001;
				8'b1001011: c <= 9'b11000001;
				8'b1101111: c <= 9'b10100111;
				8'b1101000: c <= 9'b101011101;
				8'b101100: c <= 9'b10111;
				8'b100100: c <= 9'b101101110;
				8'b1111000: c <= 9'b100000110;
				8'b1000101: c <= 9'b11111100;
				8'b1011001: c <= 9'b1111;
				8'b110100: c <= 9'b101001;
				8'b1111001: c <= 9'b111000;
				8'b1110001: c <= 9'b10111111;
				8'b1001111: c <= 9'b111011100;
				8'b1100101: c <= 9'b101111110;
				8'b1111110: c <= 9'b111001110;
				8'b1111100: c <= 9'b110011101;
				8'b1010110: c <= 9'b100001100;
				8'b110010: c <= 9'b1001111;
				8'b1101101: c <= 9'b100100010;
				8'b100011: c <= 9'b10101110;
				8'b1110101: c <= 9'b111;
				8'b1111101: c <= 9'b100101101;
				8'b101001: c <= 9'b10011011;
				8'b1010010: c <= 9'b10111101;
				8'b1011000: c <= 9'b1101111;
				8'b101110: c <= 9'b11011011;
				8'b1000001: c <= 9'b101010000;
				default: c <= 9'b0;
			endcase
			9'b1111111 : case(di)
				8'b1000011: c <= 9'b10000111;
				8'b101000: c <= 9'b111001111;
				8'b111010: c <= 9'b111101010;
				8'b110110: c <= 9'b101000010;
				8'b1100100: c <= 9'b100001;
				8'b1000000: c <= 9'b111101110;
				8'b1110110: c <= 9'b100111010;
				8'b100101: c <= 9'b101100101;
				8'b101111: c <= 9'b1001100;
				8'b100110: c <= 9'b1111001;
				8'b1100011: c <= 9'b11000100;
				8'b1001000: c <= 9'b11111011;
				8'b111000: c <= 9'b1000001;
				8'b110001: c <= 9'b100100110;
				8'b1010111: c <= 9'b1100;
				8'b1001110: c <= 9'b1000;
				8'b1101010: c <= 9'b10000011;
				8'b1001001: c <= 9'b11111001;
				8'b1100000: c <= 9'b100001001;
				8'b110111: c <= 9'b1100000;
				8'b1011101: c <= 9'b1000110;
				8'b1011011: c <= 9'b100011111;
				8'b111001: c <= 9'b101011001;
				8'b1001010: c <= 9'b110010110;
				8'b110011: c <= 9'b101110001;
				8'b1101100: c <= 9'b101010100;
				8'b1110111: c <= 9'b11010;
				8'b101011: c <= 9'b10011010;
				8'b1101011: c <= 9'b100101000;
				8'b111100: c <= 9'b110000110;
				8'b1000111: c <= 9'b1110101;
				8'b1011111: c <= 9'b100111001;
				8'b1110100: c <= 9'b1101101;
				8'b101101: c <= 9'b10000101;
				8'b1010011: c <= 9'b1110001;
				8'b1100001: c <= 9'b111110000;
				8'b110101: c <= 9'b101010;
				8'b1000100: c <= 9'b110111111;
				8'b1010001: c <= 9'b101001110;
				8'b1010100: c <= 9'b100001101;
				8'b1100110: c <= 9'b111101;
				8'b101010: c <= 9'b111111110;
				8'b1011110: c <= 9'b11100;
				8'b1100111: c <= 9'b110101111;
				8'b1011010: c <= 9'b111100110;
				8'b1000010: c <= 9'b10010110;
				8'b111101: c <= 9'b111001001;
				8'b110000: c <= 9'b100111010;
				8'b111110: c <= 9'b11101000;
				8'b1100010: c <= 9'b110100011;
				8'b1110000: c <= 9'b11100100;
				8'b1101001: c <= 9'b1100011;
				8'b1110011: c <= 9'b11010000;
				8'b1001100: c <= 9'b101110111;
				8'b100001: c <= 9'b1101111;
				8'b1000110: c <= 9'b110111;
				8'b1110010: c <= 9'b11011001;
				8'b1010000: c <= 9'b110000111;
				8'b1111010: c <= 9'b111000010;
				8'b1010101: c <= 9'b110111001;
				8'b111011: c <= 9'b111100111;
				8'b1001101: c <= 9'b11000111;
				8'b111111: c <= 9'b111010001;
				8'b1101110: c <= 9'b11000011;
				8'b1111011: c <= 9'b10;
				8'b1001011: c <= 9'b11100001;
				8'b1101111: c <= 9'b111;
				8'b1101000: c <= 9'b1000111;
				8'b101100: c <= 9'b10000000;
				8'b100100: c <= 9'b1010011;
				8'b1111000: c <= 9'b11110100;
				8'b1000101: c <= 9'b11001100;
				8'b1011001: c <= 9'b10011101;
				8'b110100: c <= 9'b11001001;
				8'b1111001: c <= 9'b111111011;
				8'b1110001: c <= 9'b11111100;
				8'b1001111: c <= 9'b100101111;
				8'b1100101: c <= 9'b110011010;
				8'b1111110: c <= 9'b111001011;
				8'b1111100: c <= 9'b1011011;
				8'b1010110: c <= 9'b111100010;
				8'b110010: c <= 9'b101111010;
				8'b1101101: c <= 9'b10011011;
				8'b100011: c <= 9'b100111110;
				8'b1110101: c <= 9'b110001011;
				8'b1111101: c <= 9'b111010111;
				8'b101001: c <= 9'b111110011;
				8'b1010010: c <= 9'b10001110;
				8'b1011000: c <= 9'b1000010;
				8'b101110: c <= 9'b11100100;
				8'b1000001: c <= 9'b11001111;
				default: c <= 9'b0;
			endcase
			9'b11110100 : case(di)
				8'b1000011: c <= 9'b110010111;
				8'b101000: c <= 9'b101110101;
				8'b111010: c <= 9'b1111100;
				8'b110110: c <= 9'b100001100;
				8'b1100100: c <= 9'b10100100;
				8'b1000000: c <= 9'b10101110;
				8'b1110110: c <= 9'b1000011;
				8'b100101: c <= 9'b111100011;
				8'b101111: c <= 9'b111001;
				8'b100110: c <= 9'b110110011;
				8'b1100011: c <= 9'b101110110;
				8'b1001000: c <= 9'b101101000;
				8'b111000: c <= 9'b1001110;
				8'b110001: c <= 9'b111100001;
				8'b1010111: c <= 9'b11100111;
				8'b1001110: c <= 9'b11001000;
				8'b1101010: c <= 9'b110010101;
				8'b1001001: c <= 9'b100110101;
				8'b1100000: c <= 9'b111011;
				8'b110111: c <= 9'b11011100;
				8'b1011101: c <= 9'b11010011;
				8'b1011011: c <= 9'b110111111;
				8'b111001: c <= 9'b1100000;
				8'b1001010: c <= 9'b101110011;
				8'b110011: c <= 9'b101010011;
				8'b1101100: c <= 9'b11110000;
				8'b1110111: c <= 9'b111100110;
				8'b101011: c <= 9'b110100;
				8'b1101011: c <= 9'b110001111;
				8'b111100: c <= 9'b110100110;
				8'b1000111: c <= 9'b10001010;
				8'b1011111: c <= 9'b110101001;
				8'b1110100: c <= 9'b100001010;
				8'b101101: c <= 9'b110000010;
				8'b1010011: c <= 9'b101000100;
				8'b1100001: c <= 9'b10110011;
				8'b110101: c <= 9'b10111100;
				8'b1000100: c <= 9'b111010110;
				8'b1010001: c <= 9'b11001101;
				8'b1010100: c <= 9'b101101010;
				8'b1100110: c <= 9'b101000011;
				8'b101010: c <= 9'b100100;
				8'b1011110: c <= 9'b1011010;
				8'b1100111: c <= 9'b111100010;
				8'b1011010: c <= 9'b110001001;
				8'b1000010: c <= 9'b101111001;
				8'b111101: c <= 9'b101101101;
				8'b110000: c <= 9'b10011011;
				8'b111110: c <= 9'b110101010;
				8'b1100010: c <= 9'b10101100;
				8'b1110000: c <= 9'b111101010;
				8'b1101001: c <= 9'b11110011;
				8'b1110011: c <= 9'b100101011;
				8'b1001100: c <= 9'b101010000;
				8'b100001: c <= 9'b100010001;
				8'b1000110: c <= 9'b10000;
				8'b1110010: c <= 9'b10101111;
				8'b1010000: c <= 9'b11001000;
				8'b1111010: c <= 9'b11010100;
				8'b1010101: c <= 9'b110110010;
				8'b111011: c <= 9'b100000111;
				8'b1001101: c <= 9'b111000010;
				8'b111111: c <= 9'b110011011;
				8'b1101110: c <= 9'b1010011;
				8'b1111011: c <= 9'b1101000;
				8'b1001011: c <= 9'b100011;
				8'b1101111: c <= 9'b1001111;
				8'b1101000: c <= 9'b10001111;
				8'b101100: c <= 9'b101111000;
				8'b100100: c <= 9'b101000110;
				8'b1111000: c <= 9'b101100000;
				8'b1000101: c <= 9'b100011001;
				8'b1011001: c <= 9'b1001000;
				8'b110100: c <= 9'b1011111;
				8'b1111001: c <= 9'b1001;
				8'b1110001: c <= 9'b110010011;
				8'b1001111: c <= 9'b110010011;
				8'b1100101: c <= 9'b110011000;
				8'b1111110: c <= 9'b110001111;
				8'b1111100: c <= 9'b10;
				8'b1010110: c <= 9'b100001111;
				8'b110010: c <= 9'b101011101;
				8'b1101101: c <= 9'b10111010;
				8'b100011: c <= 9'b1110010;
				8'b1110101: c <= 9'b1011000;
				8'b1111101: c <= 9'b1011011;
				8'b101001: c <= 9'b1111110;
				8'b1010010: c <= 9'b1000011;
				8'b1011000: c <= 9'b1000110;
				8'b101110: c <= 9'b11101001;
				8'b1000001: c <= 9'b100101101;
				default: c <= 9'b0;
			endcase
			9'b110100010 : case(di)
				8'b1000011: c <= 9'b1000011;
				8'b101000: c <= 9'b101010101;
				8'b111010: c <= 9'b101100100;
				8'b110110: c <= 9'b111010000;
				8'b1100100: c <= 9'b111100111;
				8'b1000000: c <= 9'b110110101;
				8'b1110110: c <= 9'b10010011;
				8'b100101: c <= 9'b100110101;
				8'b101111: c <= 9'b110001;
				8'b100110: c <= 9'b111111001;
				8'b1100011: c <= 9'b10111100;
				8'b1001000: c <= 9'b10100101;
				8'b111000: c <= 9'b10011111;
				8'b110001: c <= 9'b10111;
				8'b1010111: c <= 9'b10101101;
				8'b1001110: c <= 9'b10101011;
				8'b1101010: c <= 9'b100011100;
				8'b1001001: c <= 9'b10111100;
				8'b1100000: c <= 9'b100011011;
				8'b110111: c <= 9'b1110011;
				8'b1011101: c <= 9'b100100111;
				8'b1011011: c <= 9'b100011000;
				8'b111001: c <= 9'b10111000;
				8'b1001010: c <= 9'b101;
				8'b110011: c <= 9'b111111011;
				8'b1101100: c <= 9'b101100010;
				8'b1110111: c <= 9'b101001100;
				8'b101011: c <= 9'b100010100;
				8'b1101011: c <= 9'b110100001;
				8'b111100: c <= 9'b101001110;
				8'b1000111: c <= 9'b100110111;
				8'b1011111: c <= 9'b11110011;
				8'b1110100: c <= 9'b110001110;
				8'b101101: c <= 9'b111010111;
				8'b1010011: c <= 9'b10100;
				8'b1100001: c <= 9'b101011001;
				8'b110101: c <= 9'b100010010;
				8'b1000100: c <= 9'b11010111;
				8'b1010001: c <= 9'b100001011;
				8'b1010100: c <= 9'b110010;
				8'b1100110: c <= 9'b110001100;
				8'b101010: c <= 9'b11100100;
				8'b1011110: c <= 9'b10101111;
				8'b1100111: c <= 9'b10000111;
				8'b1011010: c <= 9'b101000001;
				8'b1000010: c <= 9'b110011100;
				8'b111101: c <= 9'b111100100;
				8'b110000: c <= 9'b101011010;
				8'b111110: c <= 9'b101011000;
				8'b1100010: c <= 9'b11010101;
				8'b1110000: c <= 9'b1110111;
				8'b1101001: c <= 9'b10010100;
				8'b1110011: c <= 9'b100111011;
				8'b1001100: c <= 9'b11001110;
				8'b100001: c <= 9'b101001110;
				8'b1000110: c <= 9'b1010010;
				8'b1110010: c <= 9'b100010;
				8'b1010000: c <= 9'b100010011;
				8'b1111010: c <= 9'b1111;
				8'b1010101: c <= 9'b11100000;
				8'b111011: c <= 9'b1111011;
				8'b1001101: c <= 9'b101111000;
				8'b111111: c <= 9'b110110010;
				8'b1101110: c <= 9'b11000110;
				8'b1111011: c <= 9'b100010001;
				8'b1001011: c <= 9'b1010001;
				8'b1101111: c <= 9'b101111010;
				8'b1101000: c <= 9'b101110001;
				8'b101100: c <= 9'b11110011;
				8'b100100: c <= 9'b110101101;
				8'b1111000: c <= 9'b101011101;
				8'b1000101: c <= 9'b111000011;
				8'b1011001: c <= 9'b100000111;
				8'b110100: c <= 9'b100111111;
				8'b1111001: c <= 9'b10100101;
				8'b1110001: c <= 9'b10101010;
				8'b1001111: c <= 9'b1101000;
				8'b1100101: c <= 9'b100011111;
				8'b1111110: c <= 9'b110000011;
				8'b1111100: c <= 9'b110011001;
				8'b1010110: c <= 9'b111000101;
				8'b110010: c <= 9'b110100;
				8'b1101101: c <= 9'b10111101;
				8'b100011: c <= 9'b111000011;
				8'b1110101: c <= 9'b101;
				8'b1111101: c <= 9'b1101110;
				8'b101001: c <= 9'b100010111;
				8'b1010010: c <= 9'b11000001;
				8'b1011000: c <= 9'b11101100;
				8'b101110: c <= 9'b111100111;
				8'b1000001: c <= 9'b1010101;
				default: c <= 9'b0;
			endcase
			9'b10000101 : case(di)
				8'b1000011: c <= 9'b10110010;
				8'b101000: c <= 9'b110011110;
				8'b111010: c <= 9'b100010;
				8'b110110: c <= 9'b111010111;
				8'b1100100: c <= 9'b110100010;
				8'b1000000: c <= 9'b100000101;
				8'b1110110: c <= 9'b110001100;
				8'b100101: c <= 9'b100000011;
				8'b101111: c <= 9'b111111011;
				8'b100110: c <= 9'b10000010;
				8'b1100011: c <= 9'b111010100;
				8'b1001000: c <= 9'b100001010;
				8'b111000: c <= 9'b101110000;
				8'b110001: c <= 9'b110010;
				8'b1010111: c <= 9'b10111110;
				8'b1001110: c <= 9'b110110100;
				8'b1101010: c <= 9'b10001110;
				8'b1001001: c <= 9'b100101101;
				8'b1100000: c <= 9'b110100001;
				8'b110111: c <= 9'b100000100;
				8'b1011101: c <= 9'b10000010;
				8'b1011011: c <= 9'b111110011;
				8'b111001: c <= 9'b111111010;
				8'b1001010: c <= 9'b100110;
				8'b110011: c <= 9'b100110011;
				8'b1101100: c <= 9'b1001101;
				8'b1110111: c <= 9'b110001;
				8'b101011: c <= 9'b10011011;
				8'b1101011: c <= 9'b110001001;
				8'b111100: c <= 9'b1010101;
				8'b1000111: c <= 9'b100010100;
				8'b1011111: c <= 9'b101010;
				8'b1110100: c <= 9'b11111010;
				8'b101101: c <= 9'b110110100;
				8'b1010011: c <= 9'b11111000;
				8'b1100001: c <= 9'b110001111;
				8'b110101: c <= 9'b111011111;
				8'b1000100: c <= 9'b111100010;
				8'b1010001: c <= 9'b10100011;
				8'b1010100: c <= 9'b100011001;
				8'b1100110: c <= 9'b111010010;
				8'b101010: c <= 9'b1101101;
				8'b1011110: c <= 9'b110001011;
				8'b1100111: c <= 9'b110101001;
				8'b1011010: c <= 9'b100110111;
				8'b1000010: c <= 9'b110000000;
				8'b111101: c <= 9'b101110001;
				8'b110000: c <= 9'b100001;
				8'b111110: c <= 9'b100101000;
				8'b1100010: c <= 9'b100001100;
				8'b1110000: c <= 9'b1101101;
				8'b1101001: c <= 9'b11111010;
				8'b1110011: c <= 9'b110010001;
				8'b1001100: c <= 9'b10010000;
				8'b100001: c <= 9'b101001011;
				8'b1000110: c <= 9'b1011000;
				8'b1110010: c <= 9'b1100111;
				8'b1010000: c <= 9'b10001001;
				8'b1111010: c <= 9'b101110110;
				8'b1010101: c <= 9'b110100101;
				8'b111011: c <= 9'b111111101;
				8'b1001101: c <= 9'b100000001;
				8'b111111: c <= 9'b101110110;
				8'b1101110: c <= 9'b101101110;
				8'b1111011: c <= 9'b1111001;
				8'b1001011: c <= 9'b101110100;
				8'b1101111: c <= 9'b101000111;
				8'b1101000: c <= 9'b101010001;
				8'b101100: c <= 9'b110001110;
				8'b100100: c <= 9'b110111;
				8'b1111000: c <= 9'b11110011;
				8'b1000101: c <= 9'b10100000;
				8'b1011001: c <= 9'b100100;
				8'b110100: c <= 9'b110100001;
				8'b1111001: c <= 9'b10000010;
				8'b1110001: c <= 9'b111100001;
				8'b1001111: c <= 9'b110010001;
				8'b1100101: c <= 9'b10100011;
				8'b1111110: c <= 9'b100010100;
				8'b1111100: c <= 9'b100100001;
				8'b1010110: c <= 9'b11101011;
				8'b110010: c <= 9'b111100101;
				8'b1101101: c <= 9'b101100000;
				8'b100011: c <= 9'b1000111;
				8'b1110101: c <= 9'b11010101;
				8'b1111101: c <= 9'b1001011;
				8'b101001: c <= 9'b101000001;
				8'b1010010: c <= 9'b11101011;
				8'b1011000: c <= 9'b111001100;
				8'b101110: c <= 9'b10000001;
				8'b1000001: c <= 9'b100110010;
				default: c <= 9'b0;
			endcase
			9'b101010111 : case(di)
				8'b1000011: c <= 9'b11110;
				8'b101000: c <= 9'b111111110;
				8'b111010: c <= 9'b110001100;
				8'b110110: c <= 9'b11000100;
				8'b1100100: c <= 9'b100010011;
				8'b1000000: c <= 9'b110011000;
				8'b1110110: c <= 9'b1000101;
				8'b100101: c <= 9'b110001010;
				8'b101111: c <= 9'b111101101;
				8'b100110: c <= 9'b110100100;
				8'b1100011: c <= 9'b101001011;
				8'b1001000: c <= 9'b11100111;
				8'b111000: c <= 9'b111010110;
				8'b110001: c <= 9'b110111000;
				8'b1010111: c <= 9'b110100;
				8'b1001110: c <= 9'b1110101;
				8'b1101010: c <= 9'b100;
				8'b1001001: c <= 9'b111111101;
				8'b1100000: c <= 9'b10011010;
				8'b110111: c <= 9'b101011111;
				8'b1011101: c <= 9'b100011010;
				8'b1011011: c <= 9'b10100110;
				8'b111001: c <= 9'b111100;
				8'b1001010: c <= 9'b11110101;
				8'b110011: c <= 9'b10010000;
				8'b1101100: c <= 9'b1100111;
				8'b1110111: c <= 9'b10010011;
				8'b101011: c <= 9'b111111000;
				8'b1101011: c <= 9'b101010001;
				8'b111100: c <= 9'b11111010;
				8'b1000111: c <= 9'b1111100;
				8'b1011111: c <= 9'b11101;
				8'b1110100: c <= 9'b1011111;
				8'b101101: c <= 9'b101111010;
				8'b1010011: c <= 9'b111100111;
				8'b1100001: c <= 9'b1001101;
				8'b110101: c <= 9'b1001001;
				8'b1000100: c <= 9'b11101000;
				8'b1010001: c <= 9'b10101111;
				8'b1010100: c <= 9'b1101000;
				8'b1100110: c <= 9'b111001001;
				8'b101010: c <= 9'b101010100;
				8'b1011110: c <= 9'b11001011;
				8'b1100111: c <= 9'b110000010;
				8'b1011010: c <= 9'b111011110;
				8'b1000010: c <= 9'b101000101;
				8'b111101: c <= 9'b111111010;
				8'b110000: c <= 9'b111001110;
				8'b111110: c <= 9'b11100110;
				8'b1100010: c <= 9'b111000111;
				8'b1110000: c <= 9'b110011101;
				8'b1101001: c <= 9'b10110011;
				8'b1110011: c <= 9'b11100000;
				8'b1001100: c <= 9'b1111110;
				8'b100001: c <= 9'b110000101;
				8'b1000110: c <= 9'b11010;
				8'b1110010: c <= 9'b1000000;
				8'b1010000: c <= 9'b111010111;
				8'b1111010: c <= 9'b1100011;
				8'b1010101: c <= 9'b11001001;
				8'b111011: c <= 9'b10101010;
				8'b1001101: c <= 9'b10011111;
				8'b111111: c <= 9'b110001010;
				8'b1101110: c <= 9'b11111011;
				8'b1111011: c <= 9'b100000001;
				8'b1001011: c <= 9'b111101000;
				8'b1101111: c <= 9'b101001010;
				8'b1101000: c <= 9'b100001111;
				8'b101100: c <= 9'b1101000;
				8'b100100: c <= 9'b110100001;
				8'b1111000: c <= 9'b111111110;
				8'b1000101: c <= 9'b10111011;
				8'b1011001: c <= 9'b10000101;
				8'b110100: c <= 9'b10011;
				8'b1111001: c <= 9'b10010100;
				8'b1110001: c <= 9'b1110101;
				8'b1001111: c <= 9'b101000010;
				8'b1100101: c <= 9'b1101;
				8'b1111110: c <= 9'b101100101;
				8'b1111100: c <= 9'b10110110;
				8'b1010110: c <= 9'b110100110;
				8'b110010: c <= 9'b100001111;
				8'b1101101: c <= 9'b100100010;
				8'b100011: c <= 9'b11110000;
				8'b1110101: c <= 9'b1001111;
				8'b1111101: c <= 9'b110101101;
				8'b101001: c <= 9'b1100;
				8'b1010010: c <= 9'b111110101;
				8'b1011000: c <= 9'b10000001;
				8'b101110: c <= 9'b1011011;
				8'b1000001: c <= 9'b111010111;
				default: c <= 9'b0;
			endcase
			9'b100111110 : case(di)
				8'b1000011: c <= 9'b101001110;
				8'b101000: c <= 9'b111101111;
				8'b111010: c <= 9'b111101;
				8'b110110: c <= 9'b11110111;
				8'b1100100: c <= 9'b101100000;
				8'b1000000: c <= 9'b100010001;
				8'b1110110: c <= 9'b100010111;
				8'b100101: c <= 9'b111001110;
				8'b101111: c <= 9'b100111001;
				8'b100110: c <= 9'b11111;
				8'b1100011: c <= 9'b111110101;
				8'b1001000: c <= 9'b11011;
				8'b111000: c <= 9'b110100011;
				8'b110001: c <= 9'b1000000;
				8'b1010111: c <= 9'b1001110;
				8'b1001110: c <= 9'b100100101;
				8'b1101010: c <= 9'b111110000;
				8'b1001001: c <= 9'b1001011;
				8'b1100000: c <= 9'b10010111;
				8'b110111: c <= 9'b10;
				8'b1011101: c <= 9'b1110111;
				8'b1011011: c <= 9'b11100101;
				8'b111001: c <= 9'b110000010;
				8'b1001010: c <= 9'b111010001;
				8'b110011: c <= 9'b101000011;
				8'b1101100: c <= 9'b111010000;
				8'b1110111: c <= 9'b110110000;
				8'b101011: c <= 9'b10111101;
				8'b1101011: c <= 9'b100001;
				8'b111100: c <= 9'b111111;
				8'b1000111: c <= 9'b111010100;
				8'b1011111: c <= 9'b100010101;
				8'b1110100: c <= 9'b1000001;
				8'b101101: c <= 9'b11111011;
				8'b1010011: c <= 9'b101000101;
				8'b1100001: c <= 9'b110001001;
				8'b110101: c <= 9'b110011100;
				8'b1000100: c <= 9'b111011010;
				8'b1010001: c <= 9'b10000011;
				8'b1010100: c <= 9'b1110001;
				8'b1100110: c <= 9'b101111000;
				8'b101010: c <= 9'b100001011;
				8'b1011110: c <= 9'b111111000;
				8'b1100111: c <= 9'b100011111;
				8'b1011010: c <= 9'b1001111;
				8'b1000010: c <= 9'b110101101;
				8'b111101: c <= 9'b110001110;
				8'b110000: c <= 9'b100101100;
				8'b111110: c <= 9'b1100110;
				8'b1100010: c <= 9'b100101001;
				8'b1110000: c <= 9'b110001000;
				8'b1101001: c <= 9'b11011010;
				8'b1110011: c <= 9'b111111101;
				8'b1001100: c <= 9'b10111111;
				8'b100001: c <= 9'b111100101;
				8'b1000110: c <= 9'b1011;
				8'b1110010: c <= 9'b101101010;
				8'b1010000: c <= 9'b100111;
				8'b1111010: c <= 9'b1101100;
				8'b1010101: c <= 9'b1010111;
				8'b111011: c <= 9'b110110110;
				8'b1001101: c <= 9'b1011100;
				8'b111111: c <= 9'b1110010;
				8'b1101110: c <= 9'b1101010;
				8'b1111011: c <= 9'b101001001;
				8'b1001011: c <= 9'b10110001;
				8'b1101111: c <= 9'b11001111;
				8'b1101000: c <= 9'b1001101;
				8'b101100: c <= 9'b11111010;
				8'b100100: c <= 9'b100011000;
				8'b1111000: c <= 9'b110001111;
				8'b1000101: c <= 9'b110111011;
				8'b1011001: c <= 9'b100011000;
				8'b110100: c <= 9'b100100001;
				8'b1111001: c <= 9'b101000001;
				8'b1110001: c <= 9'b10110001;
				8'b1001111: c <= 9'b10100111;
				8'b1100101: c <= 9'b10001010;
				8'b1111110: c <= 9'b11010000;
				8'b1111100: c <= 9'b110010001;
				8'b1010110: c <= 9'b11111;
				8'b110010: c <= 9'b100011001;
				8'b1101101: c <= 9'b111011111;
				8'b100011: c <= 9'b1111001;
				8'b1110101: c <= 9'b101111010;
				8'b1111101: c <= 9'b100110101;
				8'b101001: c <= 9'b10001001;
				8'b1010010: c <= 9'b111100011;
				8'b1011000: c <= 9'b111110101;
				8'b101110: c <= 9'b1111101;
				8'b1000001: c <= 9'b101000110;
				default: c <= 9'b0;
			endcase
			9'b110100000 : case(di)
				8'b1000011: c <= 9'b10100110;
				8'b101000: c <= 9'b111100110;
				8'b111010: c <= 9'b110010001;
				8'b110110: c <= 9'b110100101;
				8'b1100100: c <= 9'b11110;
				8'b1000000: c <= 9'b111110101;
				8'b1110110: c <= 9'b101101110;
				8'b100101: c <= 9'b1100000;
				8'b101111: c <= 9'b101010111;
				8'b100110: c <= 9'b10001001;
				8'b1100011: c <= 9'b11111000;
				8'b1001000: c <= 9'b10011100;
				8'b111000: c <= 9'b101101110;
				8'b110001: c <= 9'b110001110;
				8'b1010111: c <= 9'b111010000;
				8'b1001110: c <= 9'b11100000;
				8'b1101010: c <= 9'b100001001;
				8'b1001001: c <= 9'b101011101;
				8'b1100000: c <= 9'b1101001;
				8'b110111: c <= 9'b10000101;
				8'b1011101: c <= 9'b10111;
				8'b1011011: c <= 9'b1011011;
				8'b111001: c <= 9'b10011111;
				8'b1001010: c <= 9'b111110001;
				8'b110011: c <= 9'b11010011;
				8'b1101100: c <= 9'b111011110;
				8'b1110111: c <= 9'b100001001;
				8'b101011: c <= 9'b1010001;
				8'b1101011: c <= 9'b10;
				8'b111100: c <= 9'b110011011;
				8'b1000111: c <= 9'b100001011;
				8'b1011111: c <= 9'b10010011;
				8'b1110100: c <= 9'b110000010;
				8'b101101: c <= 9'b101001011;
				8'b1010011: c <= 9'b111101010;
				8'b1100001: c <= 9'b10111010;
				8'b110101: c <= 9'b10110011;
				8'b1000100: c <= 9'b110011010;
				8'b1010001: c <= 9'b111010001;
				8'b1010100: c <= 9'b111110101;
				8'b1100110: c <= 9'b10110011;
				8'b101010: c <= 9'b100110010;
				8'b1011110: c <= 9'b110000101;
				8'b1100111: c <= 9'b101101010;
				8'b1011010: c <= 9'b101110101;
				8'b1000010: c <= 9'b111100101;
				8'b111101: c <= 9'b101010;
				8'b110000: c <= 9'b111100011;
				8'b111110: c <= 9'b111100001;
				8'b1100010: c <= 9'b101011;
				8'b1110000: c <= 9'b110000010;
				8'b1101001: c <= 9'b100111101;
				8'b1110011: c <= 9'b10111110;
				8'b1001100: c <= 9'b1001100;
				8'b100001: c <= 9'b1;
				8'b1000110: c <= 9'b10100;
				8'b1110010: c <= 9'b101101110;
				8'b1010000: c <= 9'b100110101;
				8'b1111010: c <= 9'b110011000;
				8'b1010101: c <= 9'b1000101;
				8'b111011: c <= 9'b101100;
				8'b1001101: c <= 9'b11100111;
				8'b111111: c <= 9'b101100000;
				8'b1101110: c <= 9'b110000110;
				8'b1111011: c <= 9'b110000110;
				8'b1001011: c <= 9'b101011111;
				8'b1101111: c <= 9'b10101000;
				8'b1101000: c <= 9'b110010;
				8'b101100: c <= 9'b1100101;
				8'b100100: c <= 9'b100011010;
				8'b1111000: c <= 9'b111010001;
				8'b1000101: c <= 9'b100010;
				8'b1011001: c <= 9'b100101111;
				8'b110100: c <= 9'b10110011;
				8'b1111001: c <= 9'b111011011;
				8'b1110001: c <= 9'b110001001;
				8'b1001111: c <= 9'b1110001;
				8'b1100101: c <= 9'b1100100;
				8'b1111110: c <= 9'b1100;
				8'b1111100: c <= 9'b101101;
				8'b1010110: c <= 9'b111101110;
				8'b110010: c <= 9'b101010101;
				8'b1101101: c <= 9'b110010001;
				8'b100011: c <= 9'b10000011;
				8'b1110101: c <= 9'b100101000;
				8'b1111101: c <= 9'b110001010;
				8'b101001: c <= 9'b1100100;
				8'b1010010: c <= 9'b110100;
				8'b1011000: c <= 9'b110001;
				8'b101110: c <= 9'b100010101;
				8'b1000001: c <= 9'b101001010;
				default: c <= 9'b0;
			endcase
			9'b10000 : case(di)
				8'b1000011: c <= 9'b111000010;
				8'b101000: c <= 9'b110100010;
				8'b111010: c <= 9'b110100011;
				8'b110110: c <= 9'b101010000;
				8'b1100100: c <= 9'b11011101;
				8'b1000000: c <= 9'b101001111;
				8'b1110110: c <= 9'b100100011;
				8'b100101: c <= 9'b101111111;
				8'b101111: c <= 9'b111111011;
				8'b100110: c <= 9'b110101011;
				8'b1100011: c <= 9'b100100101;
				8'b1001000: c <= 9'b110000010;
				8'b111000: c <= 9'b110101010;
				8'b110001: c <= 9'b101100010;
				8'b1010111: c <= 9'b100111100;
				8'b1001110: c <= 9'b11110111;
				8'b1101010: c <= 9'b10110110;
				8'b1001001: c <= 9'b110100110;
				8'b1100000: c <= 9'b111110000;
				8'b110111: c <= 9'b111111101;
				8'b1011101: c <= 9'b10110101;
				8'b1011011: c <= 9'b100110111;
				8'b111001: c <= 9'b10001011;
				8'b1001010: c <= 9'b1100000;
				8'b110011: c <= 9'b1101110;
				8'b1101100: c <= 9'b100100010;
				8'b1110111: c <= 9'b111100010;
				8'b101011: c <= 9'b100100010;
				8'b1101011: c <= 9'b100010110;
				8'b111100: c <= 9'b1110000;
				8'b1000111: c <= 9'b111111010;
				8'b1011111: c <= 9'b110111110;
				8'b1110100: c <= 9'b1111101;
				8'b101101: c <= 9'b100010110;
				8'b1010011: c <= 9'b111010100;
				8'b1100001: c <= 9'b101111111;
				8'b110101: c <= 9'b101101001;
				8'b1000100: c <= 9'b101111001;
				8'b1010001: c <= 9'b101111000;
				8'b1010100: c <= 9'b101011;
				8'b1100110: c <= 9'b101110111;
				8'b101010: c <= 9'b11111;
				8'b1011110: c <= 9'b1001011;
				8'b1100111: c <= 9'b10000011;
				8'b1011010: c <= 9'b1010110;
				8'b1000010: c <= 9'b101011111;
				8'b111101: c <= 9'b111000010;
				8'b110000: c <= 9'b101011001;
				8'b111110: c <= 9'b1000111;
				8'b1100010: c <= 9'b10100101;
				8'b1110000: c <= 9'b1001101;
				8'b1101001: c <= 9'b110111111;
				8'b1110011: c <= 9'b100101001;
				8'b1001100: c <= 9'b110111;
				8'b100001: c <= 9'b101;
				8'b1000110: c <= 9'b111111101;
				8'b1110010: c <= 9'b1001010;
				8'b1010000: c <= 9'b101110010;
				8'b1111010: c <= 9'b111100101;
				8'b1010101: c <= 9'b100001;
				8'b111011: c <= 9'b1100000;
				8'b1001101: c <= 9'b101001011;
				8'b111111: c <= 9'b11011011;
				8'b1101110: c <= 9'b1000100;
				8'b1111011: c <= 9'b10011111;
				8'b1001011: c <= 9'b1000100;
				8'b1101111: c <= 9'b10110110;
				8'b1101000: c <= 9'b101001;
				8'b101100: c <= 9'b110000000;
				8'b100100: c <= 9'b1111010;
				8'b1111000: c <= 9'b101010100;
				8'b1000101: c <= 9'b11001000;
				8'b1011001: c <= 9'b1011100;
				8'b110100: c <= 9'b110100110;
				8'b1111001: c <= 9'b1111110;
				8'b1110001: c <= 9'b1011100;
				8'b1001111: c <= 9'b1101000;
				8'b1100101: c <= 9'b100000000;
				8'b1111110: c <= 9'b11111001;
				8'b1111100: c <= 9'b111000011;
				8'b1010110: c <= 9'b10010110;
				8'b110010: c <= 9'b11111001;
				8'b1101101: c <= 9'b110011011;
				8'b100011: c <= 9'b101101110;
				8'b1110101: c <= 9'b111001001;
				8'b1111101: c <= 9'b1100101;
				8'b101001: c <= 9'b111100000;
				8'b1010010: c <= 9'b100011010;
				8'b1011000: c <= 9'b1000011;
				8'b101110: c <= 9'b100100011;
				8'b1000001: c <= 9'b101101111;
				default: c <= 9'b0;
			endcase
			9'b101110111 : case(di)
				8'b1000011: c <= 9'b110001;
				8'b101000: c <= 9'b110001001;
				8'b111010: c <= 9'b110010111;
				8'b110110: c <= 9'b10000110;
				8'b1100100: c <= 9'b1111;
				8'b1000000: c <= 9'b100100111;
				8'b1110110: c <= 9'b111001000;
				8'b100101: c <= 9'b10010000;
				8'b101111: c <= 9'b11000100;
				8'b100110: c <= 9'b101010000;
				8'b1100011: c <= 9'b110111110;
				8'b1001000: c <= 9'b11001100;
				8'b111000: c <= 9'b11001001;
				8'b110001: c <= 9'b101010001;
				8'b1010111: c <= 9'b10010000;
				8'b1001110: c <= 9'b101010111;
				8'b1101010: c <= 9'b100100011;
				8'b1001001: c <= 9'b110111111;
				8'b1100000: c <= 9'b110010;
				8'b110111: c <= 9'b11110001;
				8'b1011101: c <= 9'b100000110;
				8'b1011011: c <= 9'b100101011;
				8'b111001: c <= 9'b1000101;
				8'b1001010: c <= 9'b11010100;
				8'b110011: c <= 9'b101000001;
				8'b1101100: c <= 9'b100101010;
				8'b1110111: c <= 9'b100010011;
				8'b101011: c <= 9'b111111;
				8'b1101011: c <= 9'b111011010;
				8'b111100: c <= 9'b10100010;
				8'b1000111: c <= 9'b11101100;
				8'b1011111: c <= 9'b1111011;
				8'b1110100: c <= 9'b110001;
				8'b101101: c <= 9'b101111001;
				8'b1010011: c <= 9'b11010;
				8'b1100001: c <= 9'b10111100;
				8'b110101: c <= 9'b1101010;
				8'b1000100: c <= 9'b100110110;
				8'b1010001: c <= 9'b10011100;
				8'b1010100: c <= 9'b11000011;
				8'b1100110: c <= 9'b111100000;
				8'b101010: c <= 9'b11100110;
				8'b1011110: c <= 9'b10111101;
				8'b1100111: c <= 9'b110111100;
				8'b1011010: c <= 9'b1101100;
				8'b1000010: c <= 9'b111001110;
				8'b111101: c <= 9'b110000101;
				8'b110000: c <= 9'b101111000;
				8'b111110: c <= 9'b1001011;
				8'b1100010: c <= 9'b111100010;
				8'b1110000: c <= 9'b111000010;
				8'b1101001: c <= 9'b111010000;
				8'b1110011: c <= 9'b100011;
				8'b1001100: c <= 9'b110110010;
				8'b100001: c <= 9'b11111101;
				8'b1000110: c <= 9'b110000011;
				8'b1110010: c <= 9'b11001110;
				8'b1010000: c <= 9'b11110001;
				8'b1111010: c <= 9'b1100100;
				8'b1010101: c <= 9'b100001111;
				8'b111011: c <= 9'b101010;
				8'b1001101: c <= 9'b111000101;
				8'b111111: c <= 9'b110011111;
				8'b1101110: c <= 9'b110011011;
				8'b1111011: c <= 9'b100100111;
				8'b1001011: c <= 9'b101100110;
				8'b1101111: c <= 9'b101111111;
				8'b1101000: c <= 9'b100010011;
				8'b101100: c <= 9'b10101111;
				8'b100100: c <= 9'b110111010;
				8'b1111000: c <= 9'b110100110;
				8'b1000101: c <= 9'b11101011;
				8'b1011001: c <= 9'b11000010;
				8'b110100: c <= 9'b110001001;
				8'b1111001: c <= 9'b10111101;
				8'b1110001: c <= 9'b101111000;
				8'b1001111: c <= 9'b1001;
				8'b1100101: c <= 9'b110101010;
				8'b1111110: c <= 9'b11110010;
				8'b1111100: c <= 9'b110110110;
				8'b1010110: c <= 9'b110100000;
				8'b110010: c <= 9'b111011100;
				8'b1101101: c <= 9'b111000011;
				8'b100011: c <= 9'b11110000;
				8'b1110101: c <= 9'b11010011;
				8'b1111101: c <= 9'b111100001;
				8'b101001: c <= 9'b110100000;
				8'b1010010: c <= 9'b101000110;
				8'b1011000: c <= 9'b110111111;
				8'b101110: c <= 9'b100101001;
				8'b1000001: c <= 9'b11000;
				default: c <= 9'b0;
			endcase
			9'b110001001 : case(di)
				8'b1000011: c <= 9'b10000101;
				8'b101000: c <= 9'b10110111;
				8'b111010: c <= 9'b11110101;
				8'b110110: c <= 9'b111101001;
				8'b1100100: c <= 9'b100000100;
				8'b1000000: c <= 9'b10010001;
				8'b1110110: c <= 9'b110000;
				8'b100101: c <= 9'b110000010;
				8'b101111: c <= 9'b110010101;
				8'b100110: c <= 9'b110100111;
				8'b1100011: c <= 9'b11100101;
				8'b1001000: c <= 9'b110001111;
				8'b111000: c <= 9'b101000100;
				8'b110001: c <= 9'b110011111;
				8'b1010111: c <= 9'b111;
				8'b1001110: c <= 9'b101110101;
				8'b1101010: c <= 9'b111000000;
				8'b1001001: c <= 9'b110101010;
				8'b1100000: c <= 9'b1111001;
				8'b110111: c <= 9'b100001010;
				8'b1011101: c <= 9'b1100011;
				8'b1011011: c <= 9'b111111;
				8'b111001: c <= 9'b111000011;
				8'b1001010: c <= 9'b101000011;
				8'b110011: c <= 9'b110100011;
				8'b1101100: c <= 9'b10000110;
				8'b1110111: c <= 9'b11001110;
				8'b101011: c <= 9'b100101111;
				8'b1101011: c <= 9'b10000;
				8'b111100: c <= 9'b110001000;
				8'b1000111: c <= 9'b11001101;
				8'b1011111: c <= 9'b10011101;
				8'b1110100: c <= 9'b101110011;
				8'b101101: c <= 9'b1111111;
				8'b1010011: c <= 9'b101100010;
				8'b1100001: c <= 9'b10011010;
				8'b110101: c <= 9'b10100100;
				8'b1000100: c <= 9'b110001100;
				8'b1010001: c <= 9'b111110000;
				8'b1010100: c <= 9'b11010001;
				8'b1100110: c <= 9'b101011110;
				8'b101010: c <= 9'b111000011;
				8'b1011110: c <= 9'b11111001;
				8'b1100111: c <= 9'b11110110;
				8'b1011010: c <= 9'b11100001;
				8'b1000010: c <= 9'b110101010;
				8'b111101: c <= 9'b100111111;
				8'b110000: c <= 9'b111000011;
				8'b111110: c <= 9'b110101010;
				8'b1100010: c <= 9'b101000100;
				8'b1110000: c <= 9'b101001010;
				8'b1101001: c <= 9'b101011000;
				8'b1110011: c <= 9'b1000001;
				8'b1001100: c <= 9'b10011111;
				8'b100001: c <= 9'b101110111;
				8'b1000110: c <= 9'b101001100;
				8'b1110010: c <= 9'b100000001;
				8'b1010000: c <= 9'b111000011;
				8'b1111010: c <= 9'b10111000;
				8'b1010101: c <= 9'b101000010;
				8'b111011: c <= 9'b10000000;
				8'b1001101: c <= 9'b11100110;
				8'b111111: c <= 9'b10110111;
				8'b1101110: c <= 9'b111101111;
				8'b1111011: c <= 9'b100011101;
				8'b1001011: c <= 9'b101001110;
				8'b1101111: c <= 9'b10111101;
				8'b1101000: c <= 9'b11010;
				8'b101100: c <= 9'b11111100;
				8'b100100: c <= 9'b110101110;
				8'b1111000: c <= 9'b11100;
				8'b1000101: c <= 9'b10101100;
				8'b1011001: c <= 9'b10101110;
				8'b110100: c <= 9'b101010;
				8'b1111001: c <= 9'b1000100;
				8'b1110001: c <= 9'b10001010;
				8'b1001111: c <= 9'b111000010;
				8'b1100101: c <= 9'b110010101;
				8'b1111110: c <= 9'b110001101;
				8'b1111100: c <= 9'b101101001;
				8'b1010110: c <= 9'b10001110;
				8'b110010: c <= 9'b1000101;
				8'b1101101: c <= 9'b110110;
				8'b100011: c <= 9'b100111100;
				8'b1110101: c <= 9'b10010110;
				8'b1111101: c <= 9'b1001100;
				8'b101001: c <= 9'b110101111;
				8'b1010010: c <= 9'b11101111;
				8'b1011000: c <= 9'b1010011;
				8'b101110: c <= 9'b100111101;
				8'b1000001: c <= 9'b110101;
				default: c <= 9'b0;
			endcase
			9'b110101111 : case(di)
				8'b1000011: c <= 9'b10110011;
				8'b101000: c <= 9'b110111111;
				8'b111010: c <= 9'b111001011;
				8'b110110: c <= 9'b111000111;
				8'b1100100: c <= 9'b110001110;
				8'b1000000: c <= 9'b10011111;
				8'b1110110: c <= 9'b110110110;
				8'b100101: c <= 9'b10110;
				8'b101111: c <= 9'b1011001;
				8'b100110: c <= 9'b100010110;
				8'b1100011: c <= 9'b1111111;
				8'b1001000: c <= 9'b1010101;
				8'b111000: c <= 9'b101001110;
				8'b110001: c <= 9'b100011011;
				8'b1010111: c <= 9'b101111111;
				8'b1001110: c <= 9'b111010001;
				8'b1101010: c <= 9'b100111110;
				8'b1001001: c <= 9'b11001101;
				8'b1100000: c <= 9'b10101110;
				8'b110111: c <= 9'b111010100;
				8'b1011101: c <= 9'b11000000;
				8'b1011011: c <= 9'b101101001;
				8'b111001: c <= 9'b11010111;
				8'b1001010: c <= 9'b100110110;
				8'b110011: c <= 9'b100101000;
				8'b1101100: c <= 9'b110100010;
				8'b1110111: c <= 9'b10001110;
				8'b101011: c <= 9'b111101111;
				8'b1101011: c <= 9'b10000110;
				8'b111100: c <= 9'b10100011;
				8'b1000111: c <= 9'b110000000;
				8'b1011111: c <= 9'b101110011;
				8'b1110100: c <= 9'b1000011;
				8'b101101: c <= 9'b110000011;
				8'b1010011: c <= 9'b10011;
				8'b1100001: c <= 9'b1001010;
				8'b110101: c <= 9'b10110011;
				8'b1000100: c <= 9'b100010011;
				8'b1010001: c <= 9'b110111111;
				8'b1010100: c <= 9'b110011;
				8'b1100110: c <= 9'b100100000;
				8'b101010: c <= 9'b111100101;
				8'b1011110: c <= 9'b110111001;
				8'b1100111: c <= 9'b100111110;
				8'b1011010: c <= 9'b11011001;
				8'b1000010: c <= 9'b100100010;
				8'b111101: c <= 9'b110001000;
				8'b110000: c <= 9'b10101111;
				8'b111110: c <= 9'b111101010;
				8'b1100010: c <= 9'b110110100;
				8'b1110000: c <= 9'b110010011;
				8'b1101001: c <= 9'b100011111;
				8'b1110011: c <= 9'b1101010;
				8'b1001100: c <= 9'b100010111;
				8'b100001: c <= 9'b11111;
				8'b1000110: c <= 9'b11111001;
				8'b1110010: c <= 9'b10000000;
				8'b1010000: c <= 9'b100010110;
				8'b1111010: c <= 9'b1100000;
				8'b1010101: c <= 9'b11000111;
				8'b111011: c <= 9'b10100010;
				8'b1001101: c <= 9'b111011011;
				8'b111111: c <= 9'b1010110;
				8'b1101110: c <= 9'b101100000;
				8'b1111011: c <= 9'b100011100;
				8'b1001011: c <= 9'b1110000;
				8'b1101111: c <= 9'b101000011;
				8'b1101000: c <= 9'b11001111;
				8'b101100: c <= 9'b10010;
				8'b100100: c <= 9'b111011111;
				8'b1111000: c <= 9'b11001100;
				8'b1000101: c <= 9'b111101;
				8'b1011001: c <= 9'b100011001;
				8'b110100: c <= 9'b1001000;
				8'b1111001: c <= 9'b100001110;
				8'b1110001: c <= 9'b11100110;
				8'b1001111: c <= 9'b100000001;
				8'b1100101: c <= 9'b10001110;
				8'b1111110: c <= 9'b1;
				8'b1111100: c <= 9'b110100100;
				8'b1010110: c <= 9'b110110111;
				8'b110010: c <= 9'b100011011;
				8'b1101101: c <= 9'b100111001;
				8'b100011: c <= 9'b10010011;
				8'b1110101: c <= 9'b111001111;
				8'b1111101: c <= 9'b100000011;
				8'b101001: c <= 9'b1000;
				8'b1010010: c <= 9'b11110000;
				8'b1011000: c <= 9'b1010101;
				8'b101110: c <= 9'b101011;
				8'b1000001: c <= 9'b11011101;
				default: c <= 9'b0;
			endcase
			9'b101110101 : case(di)
				8'b1000011: c <= 9'b1101010;
				8'b101000: c <= 9'b111001101;
				8'b111010: c <= 9'b10010101;
				8'b110110: c <= 9'b10001100;
				8'b1100100: c <= 9'b1000;
				8'b1000000: c <= 9'b10101011;
				8'b1110110: c <= 9'b110110111;
				8'b100101: c <= 9'b11110111;
				8'b101111: c <= 9'b1010101;
				8'b100110: c <= 9'b101101;
				8'b1100011: c <= 9'b11100011;
				8'b1001000: c <= 9'b11001011;
				8'b111000: c <= 9'b10110100;
				8'b110001: c <= 9'b111100000;
				8'b1010111: c <= 9'b11101000;
				8'b1001110: c <= 9'b111001011;
				8'b1101010: c <= 9'b100110010;
				8'b1001001: c <= 9'b100111011;
				8'b1100000: c <= 9'b101001110;
				8'b110111: c <= 9'b101111111;
				8'b1011101: c <= 9'b11001010;
				8'b1011011: c <= 9'b111000110;
				8'b111001: c <= 9'b100010111;
				8'b1001010: c <= 9'b111110001;
				8'b110011: c <= 9'b111011100;
				8'b1101100: c <= 9'b1100000;
				8'b1110111: c <= 9'b1010110;
				8'b101011: c <= 9'b101101101;
				8'b1101011: c <= 9'b10011000;
				8'b111100: c <= 9'b101110001;
				8'b1000111: c <= 9'b11101001;
				8'b1011111: c <= 9'b10001111;
				8'b1110100: c <= 9'b11011101;
				8'b101101: c <= 9'b111001101;
				8'b1010011: c <= 9'b10110111;
				8'b1100001: c <= 9'b100010000;
				8'b110101: c <= 9'b1000011;
				8'b1000100: c <= 9'b111100110;
				8'b1010001: c <= 9'b101001000;
				8'b1010100: c <= 9'b110100001;
				8'b1100110: c <= 9'b10110011;
				8'b101010: c <= 9'b100110110;
				8'b1011110: c <= 9'b10000001;
				8'b1100111: c <= 9'b10010;
				8'b1011010: c <= 9'b110011011;
				8'b1000010: c <= 9'b111000010;
				8'b111101: c <= 9'b1100011;
				8'b110000: c <= 9'b110100;
				8'b111110: c <= 9'b100111100;
				8'b1100010: c <= 9'b11;
				8'b1110000: c <= 9'b110111111;
				8'b1101001: c <= 9'b1011100;
				8'b1110011: c <= 9'b1100000;
				8'b1001100: c <= 9'b10110;
				8'b100001: c <= 9'b100011101;
				8'b1000110: c <= 9'b1101010;
				8'b1110010: c <= 9'b10000111;
				8'b1010000: c <= 9'b1111100;
				8'b1111010: c <= 9'b101001000;
				8'b1010101: c <= 9'b11100110;
				8'b111011: c <= 9'b111101000;
				8'b1001101: c <= 9'b1011010;
				8'b111111: c <= 9'b101001110;
				8'b1101110: c <= 9'b11001;
				8'b1111011: c <= 9'b111101110;
				8'b1001011: c <= 9'b111010111;
				8'b1101111: c <= 9'b100010011;
				8'b1101000: c <= 9'b10000101;
				8'b101100: c <= 9'b101101100;
				8'b100100: c <= 9'b100011111;
				8'b1111000: c <= 9'b11001110;
				8'b1000101: c <= 9'b111001001;
				8'b1011001: c <= 9'b100100101;
				8'b110100: c <= 9'b100111001;
				8'b1111001: c <= 9'b100111011;
				8'b1110001: c <= 9'b100001010;
				8'b1001111: c <= 9'b11011;
				8'b1100101: c <= 9'b1100110;
				8'b1111110: c <= 9'b10111001;
				8'b1111100: c <= 9'b100000011;
				8'b1010110: c <= 9'b101001;
				8'b110010: c <= 9'b101100010;
				8'b1101101: c <= 9'b101010101;
				8'b100011: c <= 9'b100100111;
				8'b1110101: c <= 9'b111001010;
				8'b1111101: c <= 9'b100100111;
				8'b101001: c <= 9'b100000011;
				8'b1010010: c <= 9'b110110110;
				8'b1011000: c <= 9'b100110;
				8'b101110: c <= 9'b1011011;
				8'b1000001: c <= 9'b1010010;
				default: c <= 9'b0;
			endcase
			9'b10101 : case(di)
				8'b1000011: c <= 9'b111001110;
				8'b101000: c <= 9'b11011001;
				8'b111010: c <= 9'b110011000;
				8'b110110: c <= 9'b11001110;
				8'b1100100: c <= 9'b100111110;
				8'b1000000: c <= 9'b111101010;
				8'b1110110: c <= 9'b111111001;
				8'b100101: c <= 9'b111000100;
				8'b101111: c <= 9'b11111100;
				8'b100110: c <= 9'b1001100;
				8'b1100011: c <= 9'b11000111;
				8'b1001000: c <= 9'b100101100;
				8'b111000: c <= 9'b100100101;
				8'b110001: c <= 9'b100110;
				8'b1010111: c <= 9'b111100101;
				8'b1001110: c <= 9'b1111000;
				8'b1101010: c <= 9'b10010000;
				8'b1001001: c <= 9'b11011101;
				8'b1100000: c <= 9'b100000101;
				8'b110111: c <= 9'b110010011;
				8'b1011101: c <= 9'b100011111;
				8'b1011011: c <= 9'b111100111;
				8'b111001: c <= 9'b110001011;
				8'b1001010: c <= 9'b101111001;
				8'b110011: c <= 9'b11110001;
				8'b1101100: c <= 9'b10101000;
				8'b1110111: c <= 9'b11001001;
				8'b101011: c <= 9'b100001111;
				8'b1101011: c <= 9'b11101100;
				8'b111100: c <= 9'b1100100;
				8'b1000111: c <= 9'b11111100;
				8'b1011111: c <= 9'b11100000;
				8'b1110100: c <= 9'b111010100;
				8'b101101: c <= 9'b10011010;
				8'b1010011: c <= 9'b1111110;
				8'b1100001: c <= 9'b100011100;
				8'b110101: c <= 9'b10111;
				8'b1000100: c <= 9'b101011011;
				8'b1010001: c <= 9'b111010010;
				8'b1010100: c <= 9'b100011010;
				8'b1100110: c <= 9'b101111111;
				8'b101010: c <= 9'b10011000;
				8'b1011110: c <= 9'b11001;
				8'b1100111: c <= 9'b101100011;
				8'b1011010: c <= 9'b101010001;
				8'b1000010: c <= 9'b100010111;
				8'b111101: c <= 9'b101111001;
				8'b110000: c <= 9'b101000001;
				8'b111110: c <= 9'b11001110;
				8'b1100010: c <= 9'b111011;
				8'b1110000: c <= 9'b101010;
				8'b1101001: c <= 9'b111100;
				8'b1110011: c <= 9'b100101000;
				8'b1001100: c <= 9'b1100;
				8'b100001: c <= 9'b11110;
				8'b1000110: c <= 9'b101100001;
				8'b1110010: c <= 9'b100100110;
				8'b1010000: c <= 9'b11100100;
				8'b1111010: c <= 9'b101001;
				8'b1010101: c <= 9'b11001110;
				8'b111011: c <= 9'b100001010;
				8'b1001101: c <= 9'b10011111;
				8'b111111: c <= 9'b111111010;
				8'b1101110: c <= 9'b101010001;
				8'b1111011: c <= 9'b101100001;
				8'b1001011: c <= 9'b110111001;
				8'b1101111: c <= 9'b100000101;
				8'b1101000: c <= 9'b101000101;
				8'b101100: c <= 9'b1011011;
				8'b100100: c <= 9'b100100;
				8'b1111000: c <= 9'b10101000;
				8'b1000101: c <= 9'b111110011;
				8'b1011001: c <= 9'b111111110;
				8'b110100: c <= 9'b10000001;
				8'b1111001: c <= 9'b10011000;
				8'b1110001: c <= 9'b110001001;
				8'b1001111: c <= 9'b111110110;
				8'b1100101: c <= 9'b101010110;
				8'b1111110: c <= 9'b111110000;
				8'b1111100: c <= 9'b100010101;
				8'b1010110: c <= 9'b100000110;
				8'b110010: c <= 9'b100110;
				8'b1101101: c <= 9'b10110001;
				8'b100011: c <= 9'b10111111;
				8'b1110101: c <= 9'b1011000;
				8'b1111101: c <= 9'b111001001;
				8'b101001: c <= 9'b1110111;
				8'b1010010: c <= 9'b11111000;
				8'b1011000: c <= 9'b1101100;
				8'b101110: c <= 9'b110101111;
				8'b1000001: c <= 9'b1110111;
				default: c <= 9'b0;
			endcase
			9'b1100011 : case(di)
				8'b1000011: c <= 9'b11000011;
				8'b101000: c <= 9'b11001001;
				8'b111010: c <= 9'b11101000;
				8'b110110: c <= 9'b11011010;
				8'b1100100: c <= 9'b101001110;
				8'b1000000: c <= 9'b111111101;
				8'b1110110: c <= 9'b1001000;
				8'b100101: c <= 9'b100011011;
				8'b101111: c <= 9'b100111110;
				8'b100110: c <= 9'b10110001;
				8'b1100011: c <= 9'b11101101;
				8'b1001000: c <= 9'b10010110;
				8'b111000: c <= 9'b1011111;
				8'b110001: c <= 9'b11001111;
				8'b1010111: c <= 9'b10110111;
				8'b1001110: c <= 9'b111100111;
				8'b1101010: c <= 9'b10101011;
				8'b1001001: c <= 9'b100111100;
				8'b1100000: c <= 9'b11001;
				8'b110111: c <= 9'b1100110;
				8'b1011101: c <= 9'b111011;
				8'b1011011: c <= 9'b110111001;
				8'b111001: c <= 9'b101010110;
				8'b1001010: c <= 9'b101100001;
				8'b110011: c <= 9'b110001000;
				8'b1101100: c <= 9'b110001110;
				8'b1110111: c <= 9'b101100100;
				8'b101011: c <= 9'b100000001;
				8'b1101011: c <= 9'b1110111;
				8'b111100: c <= 9'b10111101;
				8'b1000111: c <= 9'b101010100;
				8'b1011111: c <= 9'b11100;
				8'b1110100: c <= 9'b11010;
				8'b101101: c <= 9'b101111111;
				8'b1010011: c <= 9'b1111010;
				8'b1100001: c <= 9'b11010;
				8'b110101: c <= 9'b110111;
				8'b1000100: c <= 9'b110101111;
				8'b1010001: c <= 9'b11011011;
				8'b1010100: c <= 9'b101110111;
				8'b1100110: c <= 9'b100110111;
				8'b101010: c <= 9'b110100111;
				8'b1011110: c <= 9'b1000110;
				8'b1100111: c <= 9'b11101;
				8'b1011010: c <= 9'b11110000;
				8'b1000010: c <= 9'b100101111;
				8'b111101: c <= 9'b101011001;
				8'b110000: c <= 9'b10110110;
				8'b111110: c <= 9'b1000100;
				8'b1100010: c <= 9'b101101010;
				8'b1110000: c <= 9'b1111111;
				8'b1101001: c <= 9'b1111001;
				8'b1110011: c <= 9'b11100000;
				8'b1001100: c <= 9'b111111011;
				8'b100001: c <= 9'b11011010;
				8'b1000110: c <= 9'b1001101;
				8'b1110010: c <= 9'b110010110;
				8'b1010000: c <= 9'b1010011;
				8'b1111010: c <= 9'b101000100;
				8'b1010101: c <= 9'b110000001;
				8'b111011: c <= 9'b10100111;
				8'b1001101: c <= 9'b10001000;
				8'b111111: c <= 9'b1100101;
				8'b1101110: c <= 9'b101111110;
				8'b1111011: c <= 9'b101000100;
				8'b1001011: c <= 9'b1000001;
				8'b1101111: c <= 9'b11101000;
				8'b1101000: c <= 9'b11111011;
				8'b101100: c <= 9'b110110010;
				8'b100100: c <= 9'b101110100;
				8'b1111000: c <= 9'b111010;
				8'b1000101: c <= 9'b1000011;
				8'b1011001: c <= 9'b100010100;
				8'b110100: c <= 9'b101011010;
				8'b1111001: c <= 9'b110101101;
				8'b1110001: c <= 9'b10111001;
				8'b1001111: c <= 9'b1111111;
				8'b1100101: c <= 9'b10011001;
				8'b1111110: c <= 9'b101110110;
				8'b1111100: c <= 9'b1000001;
				8'b1010110: c <= 9'b101011010;
				8'b110010: c <= 9'b111111010;
				8'b1101101: c <= 9'b11100010;
				8'b100011: c <= 9'b110110000;
				8'b1110101: c <= 9'b10100101;
				8'b1111101: c <= 9'b101110111;
				8'b101001: c <= 9'b1110111;
				8'b1010010: c <= 9'b1100111;
				8'b1011000: c <= 9'b10110010;
				8'b101110: c <= 9'b1001010;
				8'b1000001: c <= 9'b111110011;
				default: c <= 9'b0;
			endcase
			9'b100011101 : case(di)
				8'b1000011: c <= 9'b1001110;
				8'b101000: c <= 9'b110011001;
				8'b111010: c <= 9'b101101100;
				8'b110110: c <= 9'b101001011;
				8'b1100100: c <= 9'b100101011;
				8'b1000000: c <= 9'b110100111;
				8'b1110110: c <= 9'b100000100;
				8'b100101: c <= 9'b1101;
				8'b101111: c <= 9'b111101110;
				8'b100110: c <= 9'b101101010;
				8'b1100011: c <= 9'b100110101;
				8'b1001000: c <= 9'b100001011;
				8'b111000: c <= 9'b11001000;
				8'b110001: c <= 9'b110100100;
				8'b1010111: c <= 9'b111111101;
				8'b1001110: c <= 9'b111110001;
				8'b1101010: c <= 9'b110110011;
				8'b1001001: c <= 9'b10110001;
				8'b1100000: c <= 9'b110101001;
				8'b110111: c <= 9'b111100111;
				8'b1011101: c <= 9'b110;
				8'b1011011: c <= 9'b11101101;
				8'b111001: c <= 9'b1010110;
				8'b1001010: c <= 9'b111011100;
				8'b110011: c <= 9'b11001011;
				8'b1101100: c <= 9'b111000000;
				8'b1110111: c <= 9'b100011111;
				8'b101011: c <= 9'b111101000;
				8'b1101011: c <= 9'b111111110;
				8'b111100: c <= 9'b1101;
				8'b1000111: c <= 9'b10100111;
				8'b1011111: c <= 9'b110101100;
				8'b1110100: c <= 9'b1111010;
				8'b101101: c <= 9'b110101001;
				8'b1010011: c <= 9'b110010100;
				8'b1100001: c <= 9'b101110001;
				8'b110101: c <= 9'b101101110;
				8'b1000100: c <= 9'b100101101;
				8'b1010001: c <= 9'b111001000;
				8'b1010100: c <= 9'b10000010;
				8'b1100110: c <= 9'b1001;
				8'b101010: c <= 9'b101111110;
				8'b1011110: c <= 9'b10010;
				8'b1100111: c <= 9'b111010;
				8'b1011010: c <= 9'b111001111;
				8'b1000010: c <= 9'b100100110;
				8'b111101: c <= 9'b10010111;
				8'b110000: c <= 9'b10011111;
				8'b111110: c <= 9'b111110110;
				8'b1100010: c <= 9'b10101110;
				8'b1110000: c <= 9'b101001;
				8'b1101001: c <= 9'b110100011;
				8'b1110011: c <= 9'b110110;
				8'b1001100: c <= 9'b100001;
				8'b100001: c <= 9'b101000110;
				8'b1000110: c <= 9'b111101000;
				8'b1110010: c <= 9'b110010111;
				8'b1010000: c <= 9'b110101011;
				8'b1111010: c <= 9'b10100101;
				8'b1010101: c <= 9'b100111;
				8'b111011: c <= 9'b10011100;
				8'b1001101: c <= 9'b10101000;
				8'b111111: c <= 9'b110001;
				8'b1101110: c <= 9'b111111110;
				8'b1111011: c <= 9'b101101000;
				8'b1001011: c <= 9'b1000101;
				8'b1101111: c <= 9'b11000001;
				8'b1101000: c <= 9'b110100110;
				8'b101100: c <= 9'b1110000;
				8'b100100: c <= 9'b1100100;
				8'b1111000: c <= 9'b110111010;
				8'b1000101: c <= 9'b101111010;
				8'b1011001: c <= 9'b1010011;
				8'b110100: c <= 9'b110011000;
				8'b1111001: c <= 9'b1100010;
				8'b1110001: c <= 9'b1000110;
				8'b1001111: c <= 9'b101000010;
				8'b1100101: c <= 9'b1110111;
				8'b1111110: c <= 9'b100000010;
				8'b1111100: c <= 9'b1010010;
				8'b1010110: c <= 9'b111111;
				8'b110010: c <= 9'b101101110;
				8'b1101101: c <= 9'b110011101;
				8'b100011: c <= 9'b11111001;
				8'b1110101: c <= 9'b110110111;
				8'b1111101: c <= 9'b101001010;
				8'b101001: c <= 9'b100110000;
				8'b1010010: c <= 9'b1000010;
				8'b1011000: c <= 9'b11100110;
				8'b101110: c <= 9'b110011;
				8'b1000001: c <= 9'b110001100;
				default: c <= 9'b0;
			endcase
			9'b11001011 : case(di)
				8'b1000011: c <= 9'b101111110;
				8'b101000: c <= 9'b101010101;
				8'b111010: c <= 9'b111011110;
				8'b110110: c <= 9'b1100000;
				8'b1100100: c <= 9'b101101010;
				8'b1000000: c <= 9'b11101011;
				8'b1110110: c <= 9'b111110110;
				8'b100101: c <= 9'b110011001;
				8'b101111: c <= 9'b100110100;
				8'b100110: c <= 9'b110011001;
				8'b1100011: c <= 9'b1110001;
				8'b1001000: c <= 9'b110101110;
				8'b111000: c <= 9'b1001011;
				8'b110001: c <= 9'b110010110;
				8'b1010111: c <= 9'b10011000;
				8'b1001110: c <= 9'b110111001;
				8'b1101010: c <= 9'b10111110;
				8'b1001001: c <= 9'b11010111;
				8'b1100000: c <= 9'b111111110;
				8'b110111: c <= 9'b111010000;
				8'b1011101: c <= 9'b101110100;
				8'b1011011: c <= 9'b1111010;
				8'b111001: c <= 9'b1011100;
				8'b1001010: c <= 9'b100101;
				8'b110011: c <= 9'b100111111;
				8'b1101100: c <= 9'b1100100;
				8'b1110111: c <= 9'b10110101;
				8'b101011: c <= 9'b10;
				8'b1101011: c <= 9'b111101001;
				8'b111100: c <= 9'b1100011;
				8'b1000111: c <= 9'b10110001;
				8'b1011111: c <= 9'b1001001;
				8'b1110100: c <= 9'b110101101;
				8'b101101: c <= 9'b111101000;
				8'b1010011: c <= 9'b100111100;
				8'b1100001: c <= 9'b110100000;
				8'b110101: c <= 9'b11100110;
				8'b1000100: c <= 9'b1110011;
				8'b1010001: c <= 9'b101110100;
				8'b1010100: c <= 9'b1111001;
				8'b1100110: c <= 9'b11110000;
				8'b101010: c <= 9'b101110100;
				8'b1011110: c <= 9'b110100000;
				8'b1100111: c <= 9'b1111010;
				8'b1011010: c <= 9'b111101001;
				8'b1000010: c <= 9'b11110101;
				8'b111101: c <= 9'b10111000;
				8'b110000: c <= 9'b111;
				8'b111110: c <= 9'b110001110;
				8'b1100010: c <= 9'b10011010;
				8'b1110000: c <= 9'b110110;
				8'b1101001: c <= 9'b101100010;
				8'b1110011: c <= 9'b11110011;
				8'b1001100: c <= 9'b100010100;
				8'b100001: c <= 9'b1000101;
				8'b1000110: c <= 9'b10011011;
				8'b1110010: c <= 9'b111001101;
				8'b1010000: c <= 9'b101111110;
				8'b1111010: c <= 9'b1001110;
				8'b1010101: c <= 9'b10001101;
				8'b111011: c <= 9'b1001100;
				8'b1001101: c <= 9'b1101100;
				8'b111111: c <= 9'b1000110;
				8'b1101110: c <= 9'b1001111;
				8'b1111011: c <= 9'b101101110;
				8'b1001011: c <= 9'b100110011;
				8'b1101111: c <= 9'b1001010;
				8'b1101000: c <= 9'b100110101;
				8'b101100: c <= 9'b1111001;
				8'b100100: c <= 9'b110010001;
				8'b1111000: c <= 9'b10111110;
				8'b1000101: c <= 9'b1011;
				8'b1011001: c <= 9'b100001011;
				8'b110100: c <= 9'b111110110;
				8'b1111001: c <= 9'b11000100;
				8'b1110001: c <= 9'b100001100;
				8'b1001111: c <= 9'b1001001;
				8'b1100101: c <= 9'b100001001;
				8'b1111110: c <= 9'b110100011;
				8'b1111100: c <= 9'b11110001;
				8'b1010110: c <= 9'b100000100;
				8'b110010: c <= 9'b111010100;
				8'b1101101: c <= 9'b101100101;
				8'b100011: c <= 9'b11110101;
				8'b1110101: c <= 9'b11101;
				8'b1111101: c <= 9'b100101011;
				8'b101001: c <= 9'b111000101;
				8'b1010010: c <= 9'b101011010;
				8'b1011000: c <= 9'b101110000;
				8'b101110: c <= 9'b101001010;
				8'b1000001: c <= 9'b1010111;
				default: c <= 9'b0;
			endcase
			9'b110101101 : case(di)
				8'b1000011: c <= 9'b11110000;
				8'b101000: c <= 9'b100101110;
				8'b111010: c <= 9'b110000000;
				8'b110110: c <= 9'b1001011;
				8'b1100100: c <= 9'b100111111;
				8'b1000000: c <= 9'b10111001;
				8'b1110110: c <= 9'b100111100;
				8'b100101: c <= 9'b10010100;
				8'b101111: c <= 9'b110001100;
				8'b100110: c <= 9'b11010101;
				8'b1100011: c <= 9'b100010110;
				8'b1001000: c <= 9'b100101010;
				8'b111000: c <= 9'b101000111;
				8'b110001: c <= 9'b1001100;
				8'b1010111: c <= 9'b11001000;
				8'b1001110: c <= 9'b111000011;
				8'b1101010: c <= 9'b1011111;
				8'b1001001: c <= 9'b110100101;
				8'b1100000: c <= 9'b1101101;
				8'b110111: c <= 9'b1001011;
				8'b1011101: c <= 9'b10000001;
				8'b1011011: c <= 9'b100011010;
				8'b111001: c <= 9'b101001100;
				8'b1001010: c <= 9'b111010010;
				8'b110011: c <= 9'b1001100;
				8'b1101100: c <= 9'b101001;
				8'b1110111: c <= 9'b101011110;
				8'b101011: c <= 9'b1011000;
				8'b1101011: c <= 9'b11100000;
				8'b111100: c <= 9'b1000101;
				8'b1000111: c <= 9'b10001011;
				8'b1011111: c <= 9'b110001000;
				8'b1110100: c <= 9'b1110011;
				8'b101101: c <= 9'b10010100;
				8'b1010011: c <= 9'b110100;
				8'b1100001: c <= 9'b11001111;
				8'b110101: c <= 9'b11010100;
				8'b1000100: c <= 9'b111111110;
				8'b1010001: c <= 9'b111100110;
				8'b1010100: c <= 9'b101111000;
				8'b1100110: c <= 9'b111111;
				8'b101010: c <= 9'b111001010;
				8'b1011110: c <= 9'b101001;
				8'b1100111: c <= 9'b110000001;
				8'b1011010: c <= 9'b111111110;
				8'b1000010: c <= 9'b110000001;
				8'b111101: c <= 9'b11010011;
				8'b110000: c <= 9'b101101001;
				8'b111110: c <= 9'b1000110;
				8'b1100010: c <= 9'b10110111;
				8'b1110000: c <= 9'b11001110;
				8'b1101001: c <= 9'b100110011;
				8'b1110011: c <= 9'b10010011;
				8'b1001100: c <= 9'b101111110;
				8'b100001: c <= 9'b1001110;
				8'b1000110: c <= 9'b111101101;
				8'b1110010: c <= 9'b111111110;
				8'b1010000: c <= 9'b1101111;
				8'b1111010: c <= 9'b100000001;
				8'b1010101: c <= 9'b1101110;
				8'b111011: c <= 9'b111111111;
				8'b1001101: c <= 9'b1000001;
				8'b111111: c <= 9'b110100111;
				8'b1101110: c <= 9'b111100;
				8'b1111011: c <= 9'b111011101;
				8'b1001011: c <= 9'b1001001;
				8'b1101111: c <= 9'b110011010;
				8'b1101000: c <= 9'b110101010;
				8'b101100: c <= 9'b10001000;
				8'b100100: c <= 9'b110110100;
				8'b1111000: c <= 9'b101100001;
				8'b1000101: c <= 9'b10100110;
				8'b1011001: c <= 9'b1100100;
				8'b110100: c <= 9'b110001100;
				8'b1111001: c <= 9'b10101111;
				8'b1110001: c <= 9'b10101;
				8'b1001111: c <= 9'b100110000;
				8'b1100101: c <= 9'b10011000;
				8'b1111110: c <= 9'b101110010;
				8'b1111100: c <= 9'b100110010;
				8'b1010110: c <= 9'b101101001;
				8'b110010: c <= 9'b10100100;
				8'b1101101: c <= 9'b100011010;
				8'b100011: c <= 9'b111101111;
				8'b1110101: c <= 9'b1;
				8'b1111101: c <= 9'b100111101;
				8'b101001: c <= 9'b1100000;
				8'b1010010: c <= 9'b111001001;
				8'b1011000: c <= 9'b10101000;
				8'b101110: c <= 9'b110111100;
				8'b1000001: c <= 9'b111001101;
				default: c <= 9'b0;
			endcase
			9'b110110011 : case(di)
				8'b1000011: c <= 9'b111000000;
				8'b101000: c <= 9'b111001110;
				8'b111010: c <= 9'b110100110;
				8'b110110: c <= 9'b10;
				8'b1100100: c <= 9'b110100111;
				8'b1000000: c <= 9'b11010100;
				8'b1110110: c <= 9'b100001100;
				8'b100101: c <= 9'b1100;
				8'b101111: c <= 9'b111000011;
				8'b100110: c <= 9'b111111111;
				8'b1100011: c <= 9'b100110000;
				8'b1001000: c <= 9'b111110000;
				8'b111000: c <= 9'b101111010;
				8'b110001: c <= 9'b10111000;
				8'b1010111: c <= 9'b11111101;
				8'b1001110: c <= 9'b1110101;
				8'b1101010: c <= 9'b1100011;
				8'b1001001: c <= 9'b110000011;
				8'b1100000: c <= 9'b101101110;
				8'b110111: c <= 9'b111111000;
				8'b1011101: c <= 9'b111001100;
				8'b1011011: c <= 9'b100111000;
				8'b111001: c <= 9'b10100111;
				8'b1001010: c <= 9'b111100010;
				8'b110011: c <= 9'b10111;
				8'b1101100: c <= 9'b1100001;
				8'b1110111: c <= 9'b101100;
				8'b101011: c <= 9'b100010011;
				8'b1101011: c <= 9'b10011010;
				8'b111100: c <= 9'b100111000;
				8'b1000111: c <= 9'b111011001;
				8'b1011111: c <= 9'b101000;
				8'b1110100: c <= 9'b10000101;
				8'b101101: c <= 9'b100111101;
				8'b1010011: c <= 9'b11100000;
				8'b1100001: c <= 9'b101011011;
				8'b110101: c <= 9'b100000011;
				8'b1000100: c <= 9'b100000011;
				8'b1010001: c <= 9'b111;
				8'b1010100: c <= 9'b100010;
				8'b1100110: c <= 9'b101001000;
				8'b101010: c <= 9'b10011000;
				8'b1011110: c <= 9'b10110100;
				8'b1100111: c <= 9'b110100110;
				8'b1011010: c <= 9'b1110011;
				8'b1000010: c <= 9'b101000111;
				8'b111101: c <= 9'b100101101;
				8'b110000: c <= 9'b110111111;
				8'b111110: c <= 9'b100100110;
				8'b1100010: c <= 9'b110110100;
				8'b1110000: c <= 9'b100110;
				8'b1101001: c <= 9'b101110000;
				8'b1110011: c <= 9'b11100101;
				8'b1001100: c <= 9'b110100000;
				8'b100001: c <= 9'b110110111;
				8'b1000110: c <= 9'b100111010;
				8'b1110010: c <= 9'b110111111;
				8'b1010000: c <= 9'b101001;
				8'b1111010: c <= 9'b110100011;
				8'b1010101: c <= 9'b11;
				8'b111011: c <= 9'b11101001;
				8'b1001101: c <= 9'b101011111;
				8'b111111: c <= 9'b100111011;
				8'b1101110: c <= 9'b10011100;
				8'b1111011: c <= 9'b100111011;
				8'b1001011: c <= 9'b110000110;
				8'b1101111: c <= 9'b11011100;
				8'b1101000: c <= 9'b10000;
				8'b101100: c <= 9'b111111101;
				8'b100100: c <= 9'b101100010;
				8'b1111000: c <= 9'b11000;
				8'b1000101: c <= 9'b110111111;
				8'b1011001: c <= 9'b1010010;
				8'b110100: c <= 9'b111001001;
				8'b1111001: c <= 9'b10101011;
				8'b1110001: c <= 9'b1101101;
				8'b1001111: c <= 9'b1100111;
				8'b1100101: c <= 9'b1000110;
				8'b1111110: c <= 9'b100101101;
				8'b1111100: c <= 9'b100101000;
				8'b1010110: c <= 9'b110111000;
				8'b110010: c <= 9'b111101001;
				8'b1101101: c <= 9'b111011010;
				8'b100011: c <= 9'b10111011;
				8'b1110101: c <= 9'b110100110;
				8'b1111101: c <= 9'b110000110;
				8'b101001: c <= 9'b111111000;
				8'b1010010: c <= 9'b1100010;
				8'b1011000: c <= 9'b101000100;
				8'b101110: c <= 9'b10010110;
				8'b1000001: c <= 9'b100000000;
				default: c <= 9'b0;
			endcase
			9'b101011 : case(di)
				8'b1000011: c <= 9'b101101;
				8'b101000: c <= 9'b101110100;
				8'b111010: c <= 9'b110111111;
				8'b110110: c <= 9'b111010100;
				8'b1100100: c <= 9'b101001010;
				8'b1000000: c <= 9'b101011000;
				8'b1110110: c <= 9'b111110101;
				8'b100101: c <= 9'b101010;
				8'b101111: c <= 9'b11011110;
				8'b100110: c <= 9'b100111010;
				8'b1100011: c <= 9'b1000010;
				8'b1001000: c <= 9'b111001010;
				8'b111000: c <= 9'b110010011;
				8'b110001: c <= 9'b10100101;
				8'b1010111: c <= 9'b110010110;
				8'b1001110: c <= 9'b101001010;
				8'b1101010: c <= 9'b101001000;
				8'b1001001: c <= 9'b100000101;
				8'b1100000: c <= 9'b111001100;
				8'b110111: c <= 9'b1010001;
				8'b1011101: c <= 9'b100111011;
				8'b1011011: c <= 9'b101111000;
				8'b111001: c <= 9'b111100011;
				8'b1001010: c <= 9'b110001001;
				8'b110011: c <= 9'b100001111;
				8'b1101100: c <= 9'b111000110;
				8'b1110111: c <= 9'b10100101;
				8'b101011: c <= 9'b111010010;
				8'b1101011: c <= 9'b100100;
				8'b111100: c <= 9'b111100100;
				8'b1000111: c <= 9'b110001110;
				8'b1011111: c <= 9'b10001011;
				8'b1110100: c <= 9'b10100000;
				8'b101101: c <= 9'b10111110;
				8'b1010011: c <= 9'b101010111;
				8'b1100001: c <= 9'b100011101;
				8'b110101: c <= 9'b110111001;
				8'b1000100: c <= 9'b111111011;
				8'b1010001: c <= 9'b11111010;
				8'b1010100: c <= 9'b110011;
				8'b1100110: c <= 9'b110001111;
				8'b101010: c <= 9'b110111110;
				8'b1011110: c <= 9'b100111000;
				8'b1100111: c <= 9'b101100000;
				8'b1011010: c <= 9'b100010;
				8'b1000010: c <= 9'b100001100;
				8'b111101: c <= 9'b11000;
				8'b110000: c <= 9'b100101010;
				8'b111110: c <= 9'b111010110;
				8'b1100010: c <= 9'b1000;
				8'b1110000: c <= 9'b1;
				8'b1101001: c <= 9'b110110101;
				8'b1110011: c <= 9'b1001;
				8'b1001100: c <= 9'b1011100;
				8'b100001: c <= 9'b10100101;
				8'b1000110: c <= 9'b101000101;
				8'b1110010: c <= 9'b1111101;
				8'b1010000: c <= 9'b100001;
				8'b1111010: c <= 9'b100001011;
				8'b1010101: c <= 9'b111101010;
				8'b111011: c <= 9'b11001001;
				8'b1001101: c <= 9'b110001101;
				8'b111111: c <= 9'b10100010;
				8'b1101110: c <= 9'b111111000;
				8'b1111011: c <= 9'b100110100;
				8'b1001011: c <= 9'b100101010;
				8'b1101111: c <= 9'b11011000;
				8'b1101000: c <= 9'b100000101;
				8'b101100: c <= 9'b101110101;
				8'b100100: c <= 9'b101011;
				8'b1111000: c <= 9'b100011001;
				8'b1000101: c <= 9'b1111010;
				8'b1011001: c <= 9'b101000100;
				8'b110100: c <= 9'b1000010;
				8'b1111001: c <= 9'b110111111;
				8'b1110001: c <= 9'b1010001;
				8'b1001111: c <= 9'b100101101;
				8'b1100101: c <= 9'b10011011;
				8'b1111110: c <= 9'b101000111;
				8'b1111100: c <= 9'b101101;
				8'b1010110: c <= 9'b1100001;
				8'b110010: c <= 9'b101011011;
				8'b1101101: c <= 9'b10001111;
				8'b100011: c <= 9'b110111;
				8'b1110101: c <= 9'b110111000;
				8'b1111101: c <= 9'b10001101;
				8'b101001: c <= 9'b1101010;
				8'b1010010: c <= 9'b100101;
				8'b1011000: c <= 9'b10111;
				8'b101110: c <= 9'b11101101;
				8'b1000001: c <= 9'b10101000;
				default: c <= 9'b0;
			endcase
			9'b111100110 : case(di)
				8'b1000011: c <= 9'b10001101;
				8'b101000: c <= 9'b111001001;
				8'b111010: c <= 9'b100101010;
				8'b110110: c <= 9'b10011001;
				8'b1100100: c <= 9'b111100101;
				8'b1000000: c <= 9'b1010000;
				8'b1110110: c <= 9'b1110100;
				8'b100101: c <= 9'b110111110;
				8'b101111: c <= 9'b110011001;
				8'b100110: c <= 9'b1111011;
				8'b1100011: c <= 9'b11011110;
				8'b1001000: c <= 9'b111100001;
				8'b111000: c <= 9'b111101110;
				8'b110001: c <= 9'b110101101;
				8'b1010111: c <= 9'b1111;
				8'b1001110: c <= 9'b1001001;
				8'b1101010: c <= 9'b101000011;
				8'b1001001: c <= 9'b111011111;
				8'b1100000: c <= 9'b110010001;
				8'b110111: c <= 9'b101011111;
				8'b1011101: c <= 9'b110100101;
				8'b1011011: c <= 9'b1110111;
				8'b111001: c <= 9'b10011010;
				8'b1001010: c <= 9'b100011111;
				8'b110011: c <= 9'b100011111;
				8'b1101100: c <= 9'b10100100;
				8'b1110111: c <= 9'b101100000;
				8'b101011: c <= 9'b1110001;
				8'b1101011: c <= 9'b1010110;
				8'b111100: c <= 9'b101001000;
				8'b1000111: c <= 9'b100001111;
				8'b1011111: c <= 9'b110010010;
				8'b1110100: c <= 9'b101110110;
				8'b101101: c <= 9'b10101111;
				8'b1010011: c <= 9'b111010010;
				8'b1100001: c <= 9'b11000;
				8'b110101: c <= 9'b10101000;
				8'b1000100: c <= 9'b10100;
				8'b1010001: c <= 9'b110101001;
				8'b1010100: c <= 9'b100001;
				8'b1100110: c <= 9'b10011011;
				8'b101010: c <= 9'b10111011;
				8'b1011110: c <= 9'b110011011;
				8'b1100111: c <= 9'b10001011;
				8'b1011010: c <= 9'b1011001;
				8'b1000010: c <= 9'b11011110;
				8'b111101: c <= 9'b110111110;
				8'b110000: c <= 9'b11011000;
				8'b111110: c <= 9'b1100001;
				8'b1100010: c <= 9'b11000001;
				8'b1110000: c <= 9'b11110111;
				8'b1101001: c <= 9'b111011011;
				8'b1110011: c <= 9'b10010111;
				8'b1001100: c <= 9'b11011000;
				8'b100001: c <= 9'b111111;
				8'b1000110: c <= 9'b11100100;
				8'b1110010: c <= 9'b111111;
				8'b1010000: c <= 9'b10110011;
				8'b1111010: c <= 9'b11000110;
				8'b1010101: c <= 9'b101010011;
				8'b111011: c <= 9'b101100000;
				8'b1001101: c <= 9'b10101010;
				8'b111111: c <= 9'b100011;
				8'b1101110: c <= 9'b10001110;
				8'b1111011: c <= 9'b1111110;
				8'b1001011: c <= 9'b11100001;
				8'b1101111: c <= 9'b101111000;
				8'b1101000: c <= 9'b101101100;
				8'b101100: c <= 9'b111000111;
				8'b100100: c <= 9'b11101011;
				8'b1111000: c <= 9'b10011001;
				8'b1000101: c <= 9'b101001010;
				8'b1011001: c <= 9'b100000101;
				8'b110100: c <= 9'b11101000;
				8'b1111001: c <= 9'b11011001;
				8'b1110001: c <= 9'b11001101;
				8'b1001111: c <= 9'b1011000;
				8'b1100101: c <= 9'b111100011;
				8'b1111110: c <= 9'b10000010;
				8'b1111100: c <= 9'b11011101;
				8'b1010110: c <= 9'b10010000;
				8'b110010: c <= 9'b111011101;
				8'b1101101: c <= 9'b100011010;
				8'b100011: c <= 9'b1000100;
				8'b1110101: c <= 9'b10100011;
				8'b1111101: c <= 9'b11101001;
				8'b101001: c <= 9'b10110;
				8'b1010010: c <= 9'b110100000;
				8'b1011000: c <= 9'b1111100;
				8'b101110: c <= 9'b1101111;
				8'b1000001: c <= 9'b101110100;
				default: c <= 9'b0;
			endcase
			9'b101010 : case(di)
				8'b1000011: c <= 9'b11100001;
				8'b101000: c <= 9'b1100010;
				8'b111010: c <= 9'b1110101;
				8'b110110: c <= 9'b110001111;
				8'b1100100: c <= 9'b11000;
				8'b1000000: c <= 9'b111;
				8'b1110110: c <= 9'b101010001;
				8'b100101: c <= 9'b1010010;
				8'b101111: c <= 9'b10001010;
				8'b100110: c <= 9'b111001111;
				8'b1100011: c <= 9'b100001111;
				8'b1001000: c <= 9'b10111111;
				8'b111000: c <= 9'b11101100;
				8'b110001: c <= 9'b100101110;
				8'b1010111: c <= 9'b11100;
				8'b1001110: c <= 9'b10100111;
				8'b1101010: c <= 9'b101111110;
				8'b1001001: c <= 9'b1100010;
				8'b1100000: c <= 9'b101010;
				8'b110111: c <= 9'b11100000;
				8'b1011101: c <= 9'b111000110;
				8'b1011011: c <= 9'b101010100;
				8'b111001: c <= 9'b11011000;
				8'b1001010: c <= 9'b10000110;
				8'b110011: c <= 9'b11010100;
				8'b1101100: c <= 9'b101000;
				8'b1110111: c <= 9'b101001011;
				8'b101011: c <= 9'b11011001;
				8'b1101011: c <= 9'b11100111;
				8'b111100: c <= 9'b1000001;
				8'b1000111: c <= 9'b1001;
				8'b1011111: c <= 9'b10011010;
				8'b1110100: c <= 9'b101100100;
				8'b101101: c <= 9'b110010010;
				8'b1010011: c <= 9'b101100000;
				8'b1100001: c <= 9'b11111;
				8'b110101: c <= 9'b111100;
				8'b1000100: c <= 9'b110100000;
				8'b1010001: c <= 9'b100110010;
				8'b1010100: c <= 9'b11000110;
				8'b1100110: c <= 9'b100001110;
				8'b101010: c <= 9'b10010011;
				8'b1011110: c <= 9'b10001110;
				8'b1100111: c <= 9'b11011100;
				8'b1011010: c <= 9'b1110111;
				8'b1000010: c <= 9'b111111001;
				8'b111101: c <= 9'b101011010;
				8'b110000: c <= 9'b111100010;
				8'b111110: c <= 9'b1111101;
				8'b1100010: c <= 9'b110000;
				8'b1110000: c <= 9'b110111;
				8'b1101001: c <= 9'b110011001;
				8'b1110011: c <= 9'b1;
				8'b1001100: c <= 9'b101111111;
				8'b100001: c <= 9'b11011010;
				8'b1000110: c <= 9'b10110011;
				8'b1110010: c <= 9'b11000110;
				8'b1010000: c <= 9'b1000000;
				8'b1111010: c <= 9'b10100011;
				8'b1010101: c <= 9'b1000111;
				8'b111011: c <= 9'b11101000;
				8'b1001101: c <= 9'b101011110;
				8'b111111: c <= 9'b110000111;
				8'b1101110: c <= 9'b111111001;
				8'b1111011: c <= 9'b100011111;
				8'b1001011: c <= 9'b111100010;
				8'b1101111: c <= 9'b100001101;
				8'b1101000: c <= 9'b110110101;
				8'b101100: c <= 9'b110110100;
				8'b100100: c <= 9'b1101100;
				8'b1111000: c <= 9'b10101100;
				8'b1000101: c <= 9'b111000110;
				8'b1011001: c <= 9'b100001101;
				8'b110100: c <= 9'b10101111;
				8'b1111001: c <= 9'b11010101;
				8'b1110001: c <= 9'b110000011;
				8'b1001111: c <= 9'b11000100;
				8'b1100101: c <= 9'b10010001;
				8'b1111110: c <= 9'b100110011;
				8'b1111100: c <= 9'b10010000;
				8'b1010110: c <= 9'b111100110;
				8'b110010: c <= 9'b110111010;
				8'b1101101: c <= 9'b1111000;
				8'b100011: c <= 9'b1;
				8'b1110101: c <= 9'b111010010;
				8'b1111101: c <= 9'b101001;
				8'b101001: c <= 9'b111001001;
				8'b1010010: c <= 9'b10001010;
				8'b1011000: c <= 9'b100011010;
				8'b101110: c <= 9'b111011001;
				8'b1000001: c <= 9'b101010011;
				default: c <= 9'b0;
			endcase
			9'b10001101 : case(di)
				8'b1000011: c <= 9'b1100010;
				8'b101000: c <= 9'b111100;
				8'b111010: c <= 9'b111101010;
				8'b110110: c <= 9'b11000001;
				8'b1100100: c <= 9'b11110000;
				8'b1000000: c <= 9'b111100111;
				8'b1110110: c <= 9'b110111100;
				8'b100101: c <= 9'b100101010;
				8'b101111: c <= 9'b100010010;
				8'b100110: c <= 9'b110000101;
				8'b1100011: c <= 9'b11110011;
				8'b1001000: c <= 9'b11010101;
				8'b111000: c <= 9'b1100;
				8'b110001: c <= 9'b100111000;
				8'b1010111: c <= 9'b100101010;
				8'b1001110: c <= 9'b11101000;
				8'b1101010: c <= 9'b10111011;
				8'b1001001: c <= 9'b111000010;
				8'b1100000: c <= 9'b111101001;
				8'b110111: c <= 9'b100000000;
				8'b1011101: c <= 9'b1111100;
				8'b1011011: c <= 9'b10101110;
				8'b111001: c <= 9'b11001001;
				8'b1001010: c <= 9'b110100;
				8'b110011: c <= 9'b110101111;
				8'b1101100: c <= 9'b10100111;
				8'b1110111: c <= 9'b110011110;
				8'b101011: c <= 9'b101101111;
				8'b1101011: c <= 9'b111000100;
				8'b111100: c <= 9'b101011111;
				8'b1000111: c <= 9'b101110011;
				8'b1011111: c <= 9'b101000010;
				8'b1110100: c <= 9'b101100101;
				8'b101101: c <= 9'b101011111;
				8'b1010011: c <= 9'b100110110;
				8'b1100001: c <= 9'b100010001;
				8'b110101: c <= 9'b101000111;
				8'b1000100: c <= 9'b1101110;
				8'b1010001: c <= 9'b100111111;
				8'b1010100: c <= 9'b111100;
				8'b1100110: c <= 9'b10;
				8'b101010: c <= 9'b1100100;
				8'b1011110: c <= 9'b11000;
				8'b1100111: c <= 9'b10101011;
				8'b1011010: c <= 9'b11011001;
				8'b1000010: c <= 9'b11011001;
				8'b111101: c <= 9'b10111100;
				8'b110000: c <= 9'b101011101;
				8'b111110: c <= 9'b101101010;
				8'b1100010: c <= 9'b1;
				8'b1110000: c <= 9'b10000111;
				8'b1101001: c <= 9'b111010100;
				8'b1110011: c <= 9'b101101100;
				8'b1001100: c <= 9'b10010111;
				8'b100001: c <= 9'b10111110;
				8'b1000110: c <= 9'b100110000;
				8'b1110010: c <= 9'b111011101;
				8'b1010000: c <= 9'b10001110;
				8'b1111010: c <= 9'b11111011;
				8'b1010101: c <= 9'b10100000;
				8'b111011: c <= 9'b100010011;
				8'b1001101: c <= 9'b110010101;
				8'b111111: c <= 9'b1101110;
				8'b1101110: c <= 9'b101110101;
				8'b1111011: c <= 9'b100110110;
				8'b1001011: c <= 9'b110010110;
				8'b1101111: c <= 9'b111010001;
				8'b1101000: c <= 9'b11001101;
				8'b101100: c <= 9'b1111;
				8'b100100: c <= 9'b101110001;
				8'b1111000: c <= 9'b10110;
				8'b1000101: c <= 9'b10010101;
				8'b1011001: c <= 9'b101101000;
				8'b110100: c <= 9'b1000000;
				8'b1111001: c <= 9'b10010100;
				8'b1110001: c <= 9'b11101111;
				8'b1001111: c <= 9'b111101010;
				8'b1100101: c <= 9'b1001;
				8'b1111110: c <= 9'b11110111;
				8'b1111100: c <= 9'b11111100;
				8'b1010110: c <= 9'b11000110;
				8'b110010: c <= 9'b101110100;
				8'b1101101: c <= 9'b1001001;
				8'b100011: c <= 9'b111000100;
				8'b1110101: c <= 9'b11011;
				8'b1111101: c <= 9'b110010111;
				8'b101001: c <= 9'b111111011;
				8'b1010010: c <= 9'b1101100;
				8'b1011000: c <= 9'b10111101;
				8'b101110: c <= 9'b1101110;
				8'b1000001: c <= 9'b101110101;
				default: c <= 9'b0;
			endcase
			9'b111100011 : case(di)
				8'b1000011: c <= 9'b1000110;
				8'b101000: c <= 9'b1000110;
				8'b111010: c <= 9'b10110111;
				8'b110110: c <= 9'b111000010;
				8'b1100100: c <= 9'b100000001;
				8'b1000000: c <= 9'b111100000;
				8'b1110110: c <= 9'b1001101;
				8'b100101: c <= 9'b101001;
				8'b101111: c <= 9'b111100000;
				8'b100110: c <= 9'b1101;
				8'b1100011: c <= 9'b111100010;
				8'b1001000: c <= 9'b1100100;
				8'b111000: c <= 9'b10101000;
				8'b110001: c <= 9'b110010100;
				8'b1010111: c <= 9'b11011110;
				8'b1001110: c <= 9'b101000111;
				8'b1101010: c <= 9'b111010;
				8'b1001001: c <= 9'b100000111;
				8'b1100000: c <= 9'b1000100;
				8'b110111: c <= 9'b11011011;
				8'b1011101: c <= 9'b1111000;
				8'b1011011: c <= 9'b10001101;
				8'b111001: c <= 9'b101110011;
				8'b1001010: c <= 9'b1111001;
				8'b110011: c <= 9'b1000110;
				8'b1101100: c <= 9'b110111;
				8'b1110111: c <= 9'b10110010;
				8'b101011: c <= 9'b111011100;
				8'b1101011: c <= 9'b1111;
				8'b111100: c <= 9'b100011101;
				8'b1000111: c <= 9'b111011100;
				8'b1011111: c <= 9'b11011101;
				8'b1110100: c <= 9'b101;
				8'b101101: c <= 9'b111001101;
				8'b1010011: c <= 9'b10001101;
				8'b1100001: c <= 9'b10100100;
				8'b110101: c <= 9'b11100010;
				8'b1000100: c <= 9'b100100;
				8'b1010001: c <= 9'b1001;
				8'b1010100: c <= 9'b10011000;
				8'b1100110: c <= 9'b111011;
				8'b101010: c <= 9'b1010011;
				8'b1011110: c <= 9'b1001011;
				8'b1100111: c <= 9'b1001110;
				8'b1011010: c <= 9'b11110110;
				8'b1000010: c <= 9'b111011110;
				8'b111101: c <= 9'b100011011;
				8'b110000: c <= 9'b110110010;
				8'b111110: c <= 9'b1011100;
				8'b1100010: c <= 9'b111100111;
				8'b1110000: c <= 9'b1011100;
				8'b1101001: c <= 9'b110010001;
				8'b1110011: c <= 9'b111010100;
				8'b1001100: c <= 9'b111010010;
				8'b100001: c <= 9'b110110011;
				8'b1000110: c <= 9'b101011110;
				8'b1110010: c <= 9'b1101010;
				8'b1010000: c <= 9'b111010010;
				8'b1111010: c <= 9'b1101000;
				8'b1010101: c <= 9'b10100;
				8'b111011: c <= 9'b11101101;
				8'b1001101: c <= 9'b1011000;
				8'b111111: c <= 9'b100001;
				8'b1101110: c <= 9'b1010101;
				8'b1111011: c <= 9'b110001001;
				8'b1001011: c <= 9'b11010101;
				8'b1101111: c <= 9'b110111010;
				8'b1101000: c <= 9'b1010111;
				8'b101100: c <= 9'b111110101;
				8'b100100: c <= 9'b111011111;
				8'b1111000: c <= 9'b111100000;
				8'b1000101: c <= 9'b110110011;
				8'b1011001: c <= 9'b11010011;
				8'b110100: c <= 9'b101101110;
				8'b1111001: c <= 9'b101101100;
				8'b1110001: c <= 9'b1000110;
				8'b1001111: c <= 9'b100110110;
				8'b1100101: c <= 9'b101001001;
				8'b1111110: c <= 9'b111001110;
				8'b1111100: c <= 9'b100111101;
				8'b1010110: c <= 9'b101011000;
				8'b110010: c <= 9'b100000011;
				8'b1101101: c <= 9'b100010001;
				8'b100011: c <= 9'b100011001;
				8'b1110101: c <= 9'b10010000;
				8'b1111101: c <= 9'b100110011;
				8'b101001: c <= 9'b10100100;
				8'b1010010: c <= 9'b110000001;
				8'b1011000: c <= 9'b1000000;
				8'b101110: c <= 9'b110010110;
				8'b1000001: c <= 9'b111111111;
				default: c <= 9'b0;
			endcase
			9'b100111000 : case(di)
				8'b1000011: c <= 9'b11100110;
				8'b101000: c <= 9'b110001110;
				8'b111010: c <= 9'b1110011;
				8'b110110: c <= 9'b1001110;
				8'b1100100: c <= 9'b111100000;
				8'b1000000: c <= 9'b10011011;
				8'b1110110: c <= 9'b10001101;
				8'b100101: c <= 9'b11100110;
				8'b101111: c <= 9'b101101100;
				8'b100110: c <= 9'b11011000;
				8'b1100011: c <= 9'b100011011;
				8'b1001000: c <= 9'b111110011;
				8'b111000: c <= 9'b11100010;
				8'b110001: c <= 9'b100111101;
				8'b1010111: c <= 9'b1011100;
				8'b1001110: c <= 9'b1010110;
				8'b1101010: c <= 9'b101100111;
				8'b1001001: c <= 9'b101010;
				8'b1100000: c <= 9'b110101101;
				8'b110111: c <= 9'b10001000;
				8'b1011101: c <= 9'b10110100;
				8'b1011011: c <= 9'b111000101;
				8'b111001: c <= 9'b100111;
				8'b1001010: c <= 9'b10101100;
				8'b110011: c <= 9'b10101000;
				8'b1101100: c <= 9'b100001001;
				8'b1110111: c <= 9'b110110100;
				8'b101011: c <= 9'b110110;
				8'b1101011: c <= 9'b110010101;
				8'b111100: c <= 9'b11110011;
				8'b1000111: c <= 9'b110110110;
				8'b1011111: c <= 9'b110011000;
				8'b1110100: c <= 9'b100101101;
				8'b101101: c <= 9'b100111011;
				8'b1010011: c <= 9'b110111001;
				8'b1100001: c <= 9'b101001111;
				8'b110101: c <= 9'b100001;
				8'b1000100: c <= 9'b1011010;
				8'b1010001: c <= 9'b111101010;
				8'b1010100: c <= 9'b10011101;
				8'b1100110: c <= 9'b100011010;
				8'b101010: c <= 9'b11001010;
				8'b1011110: c <= 9'b111101111;
				8'b1100111: c <= 9'b101110011;
				8'b1011010: c <= 9'b1011111;
				8'b1000010: c <= 9'b101100100;
				8'b111101: c <= 9'b100101;
				8'b110000: c <= 9'b100010110;
				8'b111110: c <= 9'b100010101;
				8'b1100010: c <= 9'b111110001;
				8'b1110000: c <= 9'b1011100;
				8'b1101001: c <= 9'b111110110;
				8'b1110011: c <= 9'b11100;
				8'b1001100: c <= 9'b100100000;
				8'b100001: c <= 9'b110;
				8'b1000110: c <= 9'b100101001;
				8'b1110010: c <= 9'b110010011;
				8'b1010000: c <= 9'b111101001;
				8'b1111010: c <= 9'b1100011;
				8'b1010101: c <= 9'b1011;
				8'b111011: c <= 9'b100011100;
				8'b1001101: c <= 9'b101011;
				8'b111111: c <= 9'b10010110;
				8'b1101110: c <= 9'b101000110;
				8'b1111011: c <= 9'b111111010;
				8'b1001011: c <= 9'b101101110;
				8'b1101111: c <= 9'b111011111;
				8'b1101000: c <= 9'b100110111;
				8'b101100: c <= 9'b11011001;
				8'b100100: c <= 9'b100000101;
				8'b1111000: c <= 9'b10011010;
				8'b1000101: c <= 9'b10101001;
				8'b1011001: c <= 9'b100111110;
				8'b110100: c <= 9'b11001010;
				8'b1111001: c <= 9'b11000;
				8'b1110001: c <= 9'b10100111;
				8'b1001111: c <= 9'b111001011;
				8'b1100101: c <= 9'b111100111;
				8'b1111110: c <= 9'b10000001;
				8'b1111100: c <= 9'b111001111;
				8'b1010110: c <= 9'b111100100;
				8'b110010: c <= 9'b100001011;
				8'b1101101: c <= 9'b100101111;
				8'b100011: c <= 9'b110110110;
				8'b1110101: c <= 9'b11011;
				8'b1111101: c <= 9'b110101100;
				8'b101001: c <= 9'b101101;
				8'b1010010: c <= 9'b1100010;
				8'b1011000: c <= 9'b10011000;
				8'b101110: c <= 9'b11000100;
				8'b1000001: c <= 9'b11100111;
				default: c <= 9'b0;
			endcase
			9'b1110000 : case(di)
				8'b1000011: c <= 9'b11001001;
				8'b101000: c <= 9'b110110100;
				8'b111010: c <= 9'b101111000;
				8'b110110: c <= 9'b101111111;
				8'b1100100: c <= 9'b111010111;
				8'b1000000: c <= 9'b110110111;
				8'b1110110: c <= 9'b11101100;
				8'b100101: c <= 9'b11101000;
				8'b101111: c <= 9'b110100000;
				8'b100110: c <= 9'b111001100;
				8'b1100011: c <= 9'b10111010;
				8'b1001000: c <= 9'b100011111;
				8'b111000: c <= 9'b1110111;
				8'b110001: c <= 9'b1101001;
				8'b1010111: c <= 9'b11100111;
				8'b1001110: c <= 9'b1011001;
				8'b1101010: c <= 9'b101000100;
				8'b1001001: c <= 9'b1011000;
				8'b1100000: c <= 9'b10001100;
				8'b110111: c <= 9'b100110101;
				8'b1011101: c <= 9'b1111000;
				8'b1011011: c <= 9'b101001011;
				8'b111001: c <= 9'b1100101;
				8'b1001010: c <= 9'b10011001;
				8'b110011: c <= 9'b110100100;
				8'b1101100: c <= 9'b11000111;
				8'b1110111: c <= 9'b101101101;
				8'b101011: c <= 9'b10111010;
				8'b1101011: c <= 9'b10101010;
				8'b111100: c <= 9'b110001000;
				8'b1000111: c <= 9'b10111110;
				8'b1011111: c <= 9'b11110100;
				8'b1110100: c <= 9'b110011101;
				8'b101101: c <= 9'b10000000;
				8'b1010011: c <= 9'b101100110;
				8'b1100001: c <= 9'b10101111;
				8'b110101: c <= 9'b100101111;
				8'b1000100: c <= 9'b100011100;
				8'b1010001: c <= 9'b11000000;
				8'b1010100: c <= 9'b101111110;
				8'b1100110: c <= 9'b11010001;
				8'b101010: c <= 9'b1110100;
				8'b1011110: c <= 9'b101100101;
				8'b1100111: c <= 9'b111001010;
				8'b1011010: c <= 9'b110100010;
				8'b1000010: c <= 9'b11100111;
				8'b111101: c <= 9'b101100001;
				8'b110000: c <= 9'b101100111;
				8'b111110: c <= 9'b1111011;
				8'b1100010: c <= 9'b101001011;
				8'b1110000: c <= 9'b101100001;
				8'b1101001: c <= 9'b11101101;
				8'b1110011: c <= 9'b1100100;
				8'b1001100: c <= 9'b1110101;
				8'b100001: c <= 9'b11001;
				8'b1000110: c <= 9'b101010010;
				8'b1110010: c <= 9'b1111110;
				8'b1010000: c <= 9'b100010111;
				8'b1111010: c <= 9'b10111110;
				8'b1010101: c <= 9'b111100001;
				8'b111011: c <= 9'b100001111;
				8'b1001101: c <= 9'b111100101;
				8'b111111: c <= 9'b101010101;
				8'b1101110: c <= 9'b111110110;
				8'b1111011: c <= 9'b1;
				8'b1001011: c <= 9'b100000101;
				8'b1101111: c <= 9'b11010111;
				8'b1101000: c <= 9'b101001011;
				8'b101100: c <= 9'b1000001;
				8'b100100: c <= 9'b1001011;
				8'b1111000: c <= 9'b100011000;
				8'b1000101: c <= 9'b11011000;
				8'b1011001: c <= 9'b100000001;
				8'b110100: c <= 9'b111111;
				8'b1111001: c <= 9'b110110010;
				8'b1110001: c <= 9'b110100;
				8'b1001111: c <= 9'b101010110;
				8'b1100101: c <= 9'b1001011;
				8'b1111110: c <= 9'b100011000;
				8'b1111100: c <= 9'b100011001;
				8'b1010110: c <= 9'b111011111;
				8'b110010: c <= 9'b111001;
				8'b1101101: c <= 9'b111100001;
				8'b100011: c <= 9'b100111011;
				8'b1110101: c <= 9'b11001010;
				8'b1111101: c <= 9'b1111;
				8'b101001: c <= 9'b101110100;
				8'b1010010: c <= 9'b111001111;
				8'b1011000: c <= 9'b11010001;
				8'b101110: c <= 9'b11011011;
				8'b1000001: c <= 9'b101111001;
				default: c <= 9'b0;
			endcase
			9'b11010010 : case(di)
				8'b1000011: c <= 9'b100110011;
				8'b101000: c <= 9'b100011000;
				8'b111010: c <= 9'b111011010;
				8'b110110: c <= 9'b101101010;
				8'b1100100: c <= 9'b111000101;
				8'b1000000: c <= 9'b111100100;
				8'b1110110: c <= 9'b111010;
				8'b100101: c <= 9'b100101100;
				8'b101111: c <= 9'b100100000;
				8'b100110: c <= 9'b1111110;
				8'b1100011: c <= 9'b10011011;
				8'b1001000: c <= 9'b10111011;
				8'b111000: c <= 9'b110111010;
				8'b110001: c <= 9'b1000101;
				8'b1010111: c <= 9'b1000000;
				8'b1001110: c <= 9'b111111011;
				8'b1101010: c <= 9'b1001011;
				8'b1001001: c <= 9'b100010010;
				8'b1100000: c <= 9'b11101101;
				8'b110111: c <= 9'b100011010;
				8'b1011101: c <= 9'b101110100;
				8'b1011011: c <= 9'b101000100;
				8'b111001: c <= 9'b110111100;
				8'b1001010: c <= 9'b1110;
				8'b110011: c <= 9'b100111001;
				8'b1101100: c <= 9'b11101001;
				8'b1110111: c <= 9'b1101001;
				8'b101011: c <= 9'b10100100;
				8'b1101011: c <= 9'b11011011;
				8'b111100: c <= 9'b100011;
				8'b1000111: c <= 9'b111001011;
				8'b1011111: c <= 9'b110101011;
				8'b1110100: c <= 9'b101111000;
				8'b101101: c <= 9'b1011010;
				8'b1010011: c <= 9'b1001011;
				8'b1100001: c <= 9'b11101101;
				8'b110101: c <= 9'b100111;
				8'b1000100: c <= 9'b11110010;
				8'b1010001: c <= 9'b101110111;
				8'b1010100: c <= 9'b101010100;
				8'b1100110: c <= 9'b110110111;
				8'b101010: c <= 9'b111011011;
				8'b1011110: c <= 9'b100001110;
				8'b1100111: c <= 9'b1011000;
				8'b1011010: c <= 9'b1000101;
				8'b1000010: c <= 9'b10011100;
				8'b111101: c <= 9'b101000001;
				8'b110000: c <= 9'b1100101;
				8'b111110: c <= 9'b1001;
				8'b1100010: c <= 9'b110101010;
				8'b1110000: c <= 9'b10001010;
				8'b1101001: c <= 9'b110010001;
				8'b1110011: c <= 9'b10001110;
				8'b1001100: c <= 9'b100111011;
				8'b100001: c <= 9'b111001101;
				8'b1000110: c <= 9'b110100001;
				8'b1110010: c <= 9'b101101000;
				8'b1010000: c <= 9'b10101100;
				8'b1111010: c <= 9'b100111;
				8'b1010101: c <= 9'b11111101;
				8'b111011: c <= 9'b11111101;
				8'b1001101: c <= 9'b1101110;
				8'b111111: c <= 9'b101110011;
				8'b1101110: c <= 9'b111010010;
				8'b1111011: c <= 9'b1101010;
				8'b1001011: c <= 9'b100000100;
				8'b1101111: c <= 9'b111011101;
				8'b1101000: c <= 9'b101100110;
				8'b101100: c <= 9'b10011100;
				8'b100100: c <= 9'b111101;
				8'b1111000: c <= 9'b111100111;
				8'b1000101: c <= 9'b101011111;
				8'b1011001: c <= 9'b1100000;
				8'b110100: c <= 9'b10000011;
				8'b1111001: c <= 9'b110000110;
				8'b1110001: c <= 9'b100110101;
				8'b1001111: c <= 9'b10101000;
				8'b1100101: c <= 9'b101110111;
				8'b1111110: c <= 9'b10001110;
				8'b1111100: c <= 9'b110100100;
				8'b1010110: c <= 9'b1001111;
				8'b110010: c <= 9'b1000111;
				8'b1101101: c <= 9'b1001000;
				8'b100011: c <= 9'b1000011;
				8'b1110101: c <= 9'b11110100;
				8'b1111101: c <= 9'b101010100;
				8'b101001: c <= 9'b100101000;
				8'b1010010: c <= 9'b10011111;
				8'b1011000: c <= 9'b1111011;
				8'b101110: c <= 9'b11110111;
				8'b1000001: c <= 9'b111100101;
				default: c <= 9'b0;
			endcase
			9'b110101001 : case(di)
				8'b1000011: c <= 9'b1011001;
				8'b101000: c <= 9'b10000110;
				8'b111010: c <= 9'b10000110;
				8'b110110: c <= 9'b100111111;
				8'b1100100: c <= 9'b1111111;
				8'b1000000: c <= 9'b10111001;
				8'b1110110: c <= 9'b11001011;
				8'b100101: c <= 9'b11111000;
				8'b101111: c <= 9'b111100000;
				8'b100110: c <= 9'b1110010;
				8'b1100011: c <= 9'b111000110;
				8'b1001000: c <= 9'b11011101;
				8'b111000: c <= 9'b100101011;
				8'b110001: c <= 9'b10111101;
				8'b1010111: c <= 9'b110100000;
				8'b1001110: c <= 9'b101010111;
				8'b1101010: c <= 9'b101011011;
				8'b1001001: c <= 9'b11101000;
				8'b1100000: c <= 9'b111010111;
				8'b110111: c <= 9'b100000110;
				8'b1011101: c <= 9'b1010011;
				8'b1011011: c <= 9'b10010001;
				8'b111001: c <= 9'b110011010;
				8'b1001010: c <= 9'b111100001;
				8'b110011: c <= 9'b100010011;
				8'b1101100: c <= 9'b11100001;
				8'b1110111: c <= 9'b1001000;
				8'b101011: c <= 9'b10111111;
				8'b1101011: c <= 9'b100111111;
				8'b111100: c <= 9'b1011000;
				8'b1000111: c <= 9'b10100110;
				8'b1011111: c <= 9'b1010110;
				8'b1110100: c <= 9'b101010001;
				8'b101101: c <= 9'b101101111;
				8'b1010011: c <= 9'b111101100;
				8'b1100001: c <= 9'b10100110;
				8'b110101: c <= 9'b10101001;
				8'b1000100: c <= 9'b101111010;
				8'b1010001: c <= 9'b110111011;
				8'b1010100: c <= 9'b1000010;
				8'b1100110: c <= 9'b110000010;
				8'b101010: c <= 9'b101101001;
				8'b1011110: c <= 9'b110;
				8'b1100111: c <= 9'b101111001;
				8'b1011010: c <= 9'b10011;
				8'b1000010: c <= 9'b100111111;
				8'b111101: c <= 9'b11100010;
				8'b110000: c <= 9'b11101100;
				8'b111110: c <= 9'b110000001;
				8'b1100010: c <= 9'b111010110;
				8'b1110000: c <= 9'b101101100;
				8'b1101001: c <= 9'b11101101;
				8'b1110011: c <= 9'b101000110;
				8'b1001100: c <= 9'b101100101;
				8'b100001: c <= 9'b110111;
				8'b1000110: c <= 9'b101010010;
				8'b1110010: c <= 9'b111110011;
				8'b1010000: c <= 9'b10110101;
				8'b1111010: c <= 9'b10011011;
				8'b1010101: c <= 9'b100111011;
				8'b111011: c <= 9'b100110100;
				8'b1001101: c <= 9'b10010100;
				8'b111111: c <= 9'b1100101;
				8'b1101110: c <= 9'b101111110;
				8'b1111011: c <= 9'b10110101;
				8'b1001011: c <= 9'b110000;
				8'b1101111: c <= 9'b110;
				8'b1101000: c <= 9'b11111011;
				8'b101100: c <= 9'b100100111;
				8'b100100: c <= 9'b1100111;
				8'b1111000: c <= 9'b110001111;
				8'b1000101: c <= 9'b11001;
				8'b1011001: c <= 9'b110000001;
				8'b110100: c <= 9'b11110101;
				8'b1111001: c <= 9'b101101001;
				8'b1110001: c <= 9'b100010011;
				8'b1001111: c <= 9'b11011110;
				8'b1100101: c <= 9'b11001001;
				8'b1111110: c <= 9'b101111110;
				8'b1111100: c <= 9'b10101011;
				8'b1010110: c <= 9'b111000101;
				8'b110010: c <= 9'b111100;
				8'b1101101: c <= 9'b111;
				8'b100011: c <= 9'b11111010;
				8'b1110101: c <= 9'b110110110;
				8'b1111101: c <= 9'b11010010;
				8'b101001: c <= 9'b10;
				8'b1010010: c <= 9'b11000010;
				8'b1011000: c <= 9'b101100101;
				8'b101110: c <= 9'b1011011;
				8'b1000001: c <= 9'b101000101;
				default: c <= 9'b0;
			endcase
			9'b1000111 : case(di)
				8'b1000011: c <= 9'b11000010;
				8'b101000: c <= 9'b111101001;
				8'b111010: c <= 9'b11111100;
				8'b110110: c <= 9'b100101000;
				8'b1100100: c <= 9'b11001100;
				8'b1000000: c <= 9'b100101100;
				8'b1110110: c <= 9'b1000001;
				8'b100101: c <= 9'b11001111;
				8'b101111: c <= 9'b100111100;
				8'b100110: c <= 9'b100111010;
				8'b1100011: c <= 9'b11;
				8'b1001000: c <= 9'b111011100;
				8'b111000: c <= 9'b10010011;
				8'b110001: c <= 9'b111100010;
				8'b1010111: c <= 9'b10011111;
				8'b1001110: c <= 9'b101011110;
				8'b1101010: c <= 9'b110101111;
				8'b1001001: c <= 9'b10001101;
				8'b1100000: c <= 9'b100001;
				8'b110111: c <= 9'b11100111;
				8'b1011101: c <= 9'b1;
				8'b1011011: c <= 9'b111101100;
				8'b111001: c <= 9'b1011000;
				8'b1001010: c <= 9'b10110101;
				8'b110011: c <= 9'b10110101;
				8'b1101100: c <= 9'b100110000;
				8'b1110111: c <= 9'b110101010;
				8'b101011: c <= 9'b101001111;
				8'b1101011: c <= 9'b10010;
				8'b111100: c <= 9'b110110110;
				8'b1000111: c <= 9'b11011011;
				8'b1011111: c <= 9'b1001101;
				8'b1110100: c <= 9'b110011110;
				8'b101101: c <= 9'b1111010;
				8'b1010011: c <= 9'b101100000;
				8'b1100001: c <= 9'b111101110;
				8'b110101: c <= 9'b100001001;
				8'b1000100: c <= 9'b10101110;
				8'b1010001: c <= 9'b10111000;
				8'b1010100: c <= 9'b1100;
				8'b1100110: c <= 9'b111111001;
				8'b101010: c <= 9'b10111111;
				8'b1011110: c <= 9'b101101010;
				8'b1100111: c <= 9'b101000010;
				8'b1011010: c <= 9'b10000001;
				8'b1000010: c <= 9'b1010010;
				8'b111101: c <= 9'b111101000;
				8'b110000: c <= 9'b101001011;
				8'b111110: c <= 9'b11111100;
				8'b1100010: c <= 9'b11100110;
				8'b1110000: c <= 9'b110100111;
				8'b1101001: c <= 9'b1010000;
				8'b1110011: c <= 9'b1111001;
				8'b1001100: c <= 9'b111100101;
				8'b100001: c <= 9'b101101111;
				8'b1000110: c <= 9'b111001;
				8'b1110010: c <= 9'b100101;
				8'b1010000: c <= 9'b1110100;
				8'b1111010: c <= 9'b11110101;
				8'b1010101: c <= 9'b100010011;
				8'b111011: c <= 9'b1011001;
				8'b1001101: c <= 9'b110110110;
				8'b111111: c <= 9'b100100110;
				8'b1101110: c <= 9'b100001100;
				8'b1111011: c <= 9'b100110101;
				8'b1001011: c <= 9'b111001001;
				8'b1101111: c <= 9'b111011010;
				8'b1101000: c <= 9'b101101010;
				8'b101100: c <= 9'b11000001;
				8'b100100: c <= 9'b11000111;
				8'b1111000: c <= 9'b10110010;
				8'b1000101: c <= 9'b110101100;
				8'b1011001: c <= 9'b111001101;
				8'b110100: c <= 9'b1001111;
				8'b1111001: c <= 9'b100001111;
				8'b1110001: c <= 9'b110001001;
				8'b1001111: c <= 9'b1110101;
				8'b1100101: c <= 9'b11100011;
				8'b1111110: c <= 9'b101100100;
				8'b1111100: c <= 9'b110000010;
				8'b1010110: c <= 9'b111101000;
				8'b110010: c <= 9'b101110010;
				8'b1101101: c <= 9'b111011001;
				8'b100011: c <= 9'b11100000;
				8'b1110101: c <= 9'b110011111;
				8'b1111101: c <= 9'b1111101;
				8'b101001: c <= 9'b11001100;
				8'b1010010: c <= 9'b101100;
				8'b1011000: c <= 9'b10110011;
				8'b101110: c <= 9'b11100001;
				8'b1000001: c <= 9'b11111;
				default: c <= 9'b0;
			endcase
			9'b101100011 : case(di)
				8'b1000011: c <= 9'b1100111;
				8'b101000: c <= 9'b11100100;
				8'b111010: c <= 9'b101010100;
				8'b110110: c <= 9'b100010010;
				8'b1100100: c <= 9'b10001101;
				8'b1000000: c <= 9'b11000;
				8'b1110110: c <= 9'b101011111;
				8'b100101: c <= 9'b10111101;
				8'b101111: c <= 9'b100100110;
				8'b100110: c <= 9'b111000;
				8'b1100011: c <= 9'b11101001;
				8'b1001000: c <= 9'b1001101;
				8'b111000: c <= 9'b1111101;
				8'b110001: c <= 9'b111101010;
				8'b1010111: c <= 9'b1001111;
				8'b1001110: c <= 9'b101101101;
				8'b1101010: c <= 9'b110;
				8'b1001001: c <= 9'b100001111;
				8'b1100000: c <= 9'b100001001;
				8'b110111: c <= 9'b101111010;
				8'b1011101: c <= 9'b101011110;
				8'b1011011: c <= 9'b1101110;
				8'b111001: c <= 9'b11110110;
				8'b1001010: c <= 9'b111011100;
				8'b110011: c <= 9'b110101001;
				8'b1101100: c <= 9'b111001100;
				8'b1110111: c <= 9'b10110011;
				8'b101011: c <= 9'b110100100;
				8'b1101011: c <= 9'b11000001;
				8'b111100: c <= 9'b100101101;
				8'b1000111: c <= 9'b10000111;
				8'b1011111: c <= 9'b100111100;
				8'b1110100: c <= 9'b110111110;
				8'b101101: c <= 9'b111100001;
				8'b1010011: c <= 9'b10011001;
				8'b1100001: c <= 9'b101100100;
				8'b110101: c <= 9'b1000001;
				8'b1000100: c <= 9'b10010;
				8'b1010001: c <= 9'b100001101;
				8'b1010100: c <= 9'b11001110;
				8'b1100110: c <= 9'b1100;
				8'b101010: c <= 9'b11111101;
				8'b1011110: c <= 9'b100000101;
				8'b1100111: c <= 9'b111010001;
				8'b1011010: c <= 9'b111110000;
				8'b1000010: c <= 9'b10110;
				8'b111101: c <= 9'b110111111;
				8'b110000: c <= 9'b1101000;
				8'b111110: c <= 9'b11011011;
				8'b1100010: c <= 9'b101001111;
				8'b1110000: c <= 9'b11011101;
				8'b1101001: c <= 9'b101110101;
				8'b1110011: c <= 9'b110010100;
				8'b1001100: c <= 9'b110000111;
				8'b100001: c <= 9'b10110011;
				8'b1000110: c <= 9'b100011100;
				8'b1110010: c <= 9'b10010110;
				8'b1010000: c <= 9'b11100011;
				8'b1111010: c <= 9'b1100010;
				8'b1010101: c <= 9'b1011001;
				8'b111011: c <= 9'b11111010;
				8'b1001101: c <= 9'b1001011;
				8'b111111: c <= 9'b111010001;
				8'b1101110: c <= 9'b100110000;
				8'b1111011: c <= 9'b111111101;
				8'b1001011: c <= 9'b1100111;
				8'b1101111: c <= 9'b10110001;
				8'b1101000: c <= 9'b101110000;
				8'b101100: c <= 9'b101001111;
				8'b100100: c <= 9'b10000110;
				8'b1111000: c <= 9'b100101010;
				8'b1000101: c <= 9'b101010110;
				8'b1011001: c <= 9'b100010110;
				8'b110100: c <= 9'b10010110;
				8'b1111001: c <= 9'b10001100;
				8'b1110001: c <= 9'b100100000;
				8'b1001111: c <= 9'b11110011;
				8'b1100101: c <= 9'b11110001;
				8'b1111110: c <= 9'b1011111;
				8'b1111100: c <= 9'b11011100;
				8'b1010110: c <= 9'b10001110;
				8'b110010: c <= 9'b110111001;
				8'b1101101: c <= 9'b111101100;
				8'b100011: c <= 9'b101100010;
				8'b1110101: c <= 9'b11100000;
				8'b1111101: c <= 9'b1111;
				8'b101001: c <= 9'b111100011;
				8'b1010010: c <= 9'b101100;
				8'b1011000: c <= 9'b111001110;
				8'b101110: c <= 9'b100011100;
				8'b1000001: c <= 9'b11110100;
				default: c <= 9'b0;
			endcase
			9'b111110101 : case(di)
				8'b1000011: c <= 9'b100101001;
				8'b101000: c <= 9'b1110;
				8'b111010: c <= 9'b1001;
				8'b110110: c <= 9'b10010001;
				8'b1100100: c <= 9'b110100000;
				8'b1000000: c <= 9'b101000011;
				8'b1110110: c <= 9'b1000111;
				8'b100101: c <= 9'b1011010;
				8'b101111: c <= 9'b1001111;
				8'b100110: c <= 9'b101001111;
				8'b1100011: c <= 9'b10110111;
				8'b1001000: c <= 9'b10101110;
				8'b111000: c <= 9'b1110010;
				8'b110001: c <= 9'b11011001;
				8'b1010111: c <= 9'b10101101;
				8'b1001110: c <= 9'b100010001;
				8'b1101010: c <= 9'b11000111;
				8'b1001001: c <= 9'b11010011;
				8'b1100000: c <= 9'b110100100;
				8'b110111: c <= 9'b10101110;
				8'b1011101: c <= 9'b10101100;
				8'b1011011: c <= 9'b111111011;
				8'b111001: c <= 9'b10100010;
				8'b1001010: c <= 9'b110100;
				8'b110011: c <= 9'b10110;
				8'b1101100: c <= 9'b110000010;
				8'b1110111: c <= 9'b10010;
				8'b101011: c <= 9'b10101100;
				8'b1101011: c <= 9'b111000100;
				8'b111100: c <= 9'b10100;
				8'b1000111: c <= 9'b11110101;
				8'b1011111: c <= 9'b101110100;
				8'b1110100: c <= 9'b1101;
				8'b101101: c <= 9'b111111111;
				8'b1010011: c <= 9'b101110101;
				8'b1100001: c <= 9'b11100;
				8'b110101: c <= 9'b1110101;
				8'b1000100: c <= 9'b100111101;
				8'b1010001: c <= 9'b101100110;
				8'b1010100: c <= 9'b110100;
				8'b1100110: c <= 9'b1011100;
				8'b101010: c <= 9'b100011010;
				8'b1011110: c <= 9'b11101011;
				8'b1100111: c <= 9'b100010001;
				8'b1011010: c <= 9'b110100110;
				8'b1000010: c <= 9'b100011010;
				8'b111101: c <= 9'b100111;
				8'b110000: c <= 9'b11101111;
				8'b111110: c <= 9'b1101101;
				8'b1100010: c <= 9'b1010010;
				8'b1110000: c <= 9'b111011111;
				8'b1101001: c <= 9'b100010110;
				8'b1110011: c <= 9'b100000000;
				8'b1001100: c <= 9'b111011101;
				8'b100001: c <= 9'b11011101;
				8'b1000110: c <= 9'b10001111;
				8'b1110010: c <= 9'b111011011;
				8'b1010000: c <= 9'b110010100;
				8'b1111010: c <= 9'b101110010;
				8'b1010101: c <= 9'b111101100;
				8'b111011: c <= 9'b100111000;
				8'b1001101: c <= 9'b1111000;
				8'b111111: c <= 9'b100000111;
				8'b1101110: c <= 9'b111000101;
				8'b1111011: c <= 9'b1101110;
				8'b1001011: c <= 9'b110100000;
				8'b1101111: c <= 9'b10;
				8'b1101000: c <= 9'b101000100;
				8'b101100: c <= 9'b101001010;
				8'b100100: c <= 9'b110001011;
				8'b1111000: c <= 9'b10100010;
				8'b1000101: c <= 9'b100010101;
				8'b1011001: c <= 9'b11101100;
				8'b110100: c <= 9'b100100011;
				8'b1111001: c <= 9'b1010110;
				8'b1110001: c <= 9'b11011010;
				8'b1001111: c <= 9'b1101110;
				8'b1100101: c <= 9'b100100;
				8'b1111110: c <= 9'b100111101;
				8'b1111100: c <= 9'b111100110;
				8'b1010110: c <= 9'b1000;
				8'b110010: c <= 9'b1110101;
				8'b1101101: c <= 9'b1101110;
				8'b100011: c <= 9'b1111000;
				8'b1110101: c <= 9'b111000101;
				8'b1111101: c <= 9'b10101111;
				8'b101001: c <= 9'b101110111;
				8'b1010010: c <= 9'b1111111;
				8'b1011000: c <= 9'b110011;
				8'b101110: c <= 9'b10000;
				8'b1000001: c <= 9'b1011100;
				default: c <= 9'b0;
			endcase
			9'b1000001 : case(di)
				8'b1000011: c <= 9'b111100010;
				8'b101000: c <= 9'b100010001;
				8'b111010: c <= 9'b10100011;
				8'b110110: c <= 9'b11110110;
				8'b1100100: c <= 9'b1001101;
				8'b1000000: c <= 9'b111111;
				8'b1110110: c <= 9'b1000001;
				8'b100101: c <= 9'b1001110;
				8'b101111: c <= 9'b11001010;
				8'b100110: c <= 9'b11100010;
				8'b1100011: c <= 9'b11011110;
				8'b1001000: c <= 9'b100110101;
				8'b111000: c <= 9'b11110111;
				8'b110001: c <= 9'b101111111;
				8'b1010111: c <= 9'b100000001;
				8'b1001110: c <= 9'b111100000;
				8'b1101010: c <= 9'b1010000;
				8'b1001001: c <= 9'b1000;
				8'b1100000: c <= 9'b110011;
				8'b110111: c <= 9'b1010010;
				8'b1011101: c <= 9'b100101011;
				8'b1011011: c <= 9'b10010001;
				8'b111001: c <= 9'b10101011;
				8'b1001010: c <= 9'b110001110;
				8'b110011: c <= 9'b101010;
				8'b1101100: c <= 9'b111110011;
				8'b1110111: c <= 9'b100101;
				8'b101011: c <= 9'b111011110;
				8'b1101011: c <= 9'b1110000;
				8'b111100: c <= 9'b100111010;
				8'b1000111: c <= 9'b10001101;
				8'b1011111: c <= 9'b110110;
				8'b1110100: c <= 9'b100100;
				8'b101101: c <= 9'b10100;
				8'b1010011: c <= 9'b100010111;
				8'b1100001: c <= 9'b100100011;
				8'b110101: c <= 9'b110001100;
				8'b1000100: c <= 9'b10001011;
				8'b1010001: c <= 9'b111110001;
				8'b1010100: c <= 9'b101001010;
				8'b1100110: c <= 9'b1001011;
				8'b101010: c <= 9'b10101111;
				8'b1011110: c <= 9'b10011100;
				8'b1100111: c <= 9'b11000001;
				8'b1011010: c <= 9'b100100000;
				8'b1000010: c <= 9'b110110111;
				8'b111101: c <= 9'b10100100;
				8'b110000: c <= 9'b11100010;
				8'b111110: c <= 9'b10011;
				8'b1100010: c <= 9'b1110011;
				8'b1110000: c <= 9'b1011100;
				8'b1101001: c <= 9'b101011101;
				8'b1110011: c <= 9'b110000110;
				8'b1001100: c <= 9'b111001011;
				8'b100001: c <= 9'b101001;
				8'b1000110: c <= 9'b110010010;
				8'b1110010: c <= 9'b111101000;
				8'b1010000: c <= 9'b100001100;
				8'b1111010: c <= 9'b1100010;
				8'b1010101: c <= 9'b110111011;
				8'b111011: c <= 9'b10010011;
				8'b1001101: c <= 9'b111111110;
				8'b111111: c <= 9'b111110001;
				8'b1101110: c <= 9'b110110101;
				8'b1111011: c <= 9'b100101110;
				8'b1001011: c <= 9'b10110011;
				8'b1101111: c <= 9'b101011111;
				8'b1101000: c <= 9'b111110101;
				8'b101100: c <= 9'b1000010;
				8'b100100: c <= 9'b110101110;
				8'b1111000: c <= 9'b101101;
				8'b1000101: c <= 9'b1111110;
				8'b1011001: c <= 9'b11111011;
				8'b110100: c <= 9'b1;
				8'b1111001: c <= 9'b101101111;
				8'b1110001: c <= 9'b101110011;
				8'b1001111: c <= 9'b100000010;
				8'b1100101: c <= 9'b1001011;
				8'b1111110: c <= 9'b10011100;
				8'b1111100: c <= 9'b110001011;
				8'b1010110: c <= 9'b110110111;
				8'b110010: c <= 9'b10111100;
				8'b1101101: c <= 9'b110011010;
				8'b100011: c <= 9'b110010110;
				8'b1110101: c <= 9'b11;
				8'b1111101: c <= 9'b10110011;
				8'b101001: c <= 9'b1101111;
				8'b1010010: c <= 9'b1100101;
				8'b1011000: c <= 9'b111001001;
				8'b101110: c <= 9'b10110010;
				8'b1000001: c <= 9'b10111001;
				default: c <= 9'b0;
			endcase
			9'b110000111 : case(di)
				8'b1000011: c <= 9'b110100110;
				8'b101000: c <= 9'b11100100;
				8'b111010: c <= 9'b1011011;
				8'b110110: c <= 9'b1011;
				8'b1100100: c <= 9'b1001000;
				8'b1000000: c <= 9'b11110000;
				8'b1110110: c <= 9'b110111000;
				8'b100101: c <= 9'b101010110;
				8'b101111: c <= 9'b1010000;
				8'b100110: c <= 9'b11101000;
				8'b1100011: c <= 9'b110000011;
				8'b1001000: c <= 9'b11010000;
				8'b111000: c <= 9'b100011111;
				8'b110001: c <= 9'b111011110;
				8'b1010111: c <= 9'b110100001;
				8'b1001110: c <= 9'b1100111;
				8'b1101010: c <= 9'b111010100;
				8'b1001001: c <= 9'b1111100;
				8'b1100000: c <= 9'b1011100;
				8'b110111: c <= 9'b111001101;
				8'b1011101: c <= 9'b1010111;
				8'b1011011: c <= 9'b100101000;
				8'b111001: c <= 9'b101001111;
				8'b1001010: c <= 9'b101000110;
				8'b110011: c <= 9'b111011001;
				8'b1101100: c <= 9'b100010110;
				8'b1110111: c <= 9'b110111;
				8'b101011: c <= 9'b10101101;
				8'b1101011: c <= 9'b110100111;
				8'b111100: c <= 9'b111101101;
				8'b1000111: c <= 9'b111010111;
				8'b1011111: c <= 9'b1011011;
				8'b1110100: c <= 9'b1111;
				8'b101101: c <= 9'b11101101;
				8'b1010011: c <= 9'b10101001;
				8'b1100001: c <= 9'b110110101;
				8'b110101: c <= 9'b1011011;
				8'b1000100: c <= 9'b110110011;
				8'b1010001: c <= 9'b111101111;
				8'b1010100: c <= 9'b1110000;
				8'b1100110: c <= 9'b110001000;
				8'b101010: c <= 9'b1000011;
				8'b1011110: c <= 9'b101110000;
				8'b1100111: c <= 9'b111111011;
				8'b1011010: c <= 9'b11100001;
				8'b1000010: c <= 9'b10111011;
				8'b111101: c <= 9'b1001;
				8'b110000: c <= 9'b110011110;
				8'b111110: c <= 9'b11111;
				8'b1100010: c <= 9'b11101;
				8'b1110000: c <= 9'b11;
				8'b1101001: c <= 9'b110101100;
				8'b1110011: c <= 9'b1010101;
				8'b1001100: c <= 9'b110111010;
				8'b100001: c <= 9'b10010111;
				8'b1000110: c <= 9'b110010110;
				8'b1110010: c <= 9'b110000101;
				8'b1010000: c <= 9'b101110101;
				8'b1111010: c <= 9'b101011111;
				8'b1010101: c <= 9'b10000010;
				8'b111011: c <= 9'b110001100;
				8'b1001101: c <= 9'b10110011;
				8'b111111: c <= 9'b11010101;
				8'b1101110: c <= 9'b101101010;
				8'b1111011: c <= 9'b101110000;
				8'b1001011: c <= 9'b101001;
				8'b1101111: c <= 9'b101011;
				8'b1101000: c <= 9'b10111111;
				8'b101100: c <= 9'b101111110;
				8'b100100: c <= 9'b110011110;
				8'b1111000: c <= 9'b11001000;
				8'b1000101: c <= 9'b10001010;
				8'b1011001: c <= 9'b10010;
				8'b110100: c <= 9'b110101100;
				8'b1111001: c <= 9'b11100010;
				8'b1110001: c <= 9'b1001000;
				8'b1001111: c <= 9'b10110110;
				8'b1100101: c <= 9'b110100110;
				8'b1111110: c <= 9'b10000111;
				8'b1111100: c <= 9'b10101;
				8'b1010110: c <= 9'b100110100;
				8'b110010: c <= 9'b10110011;
				8'b1101101: c <= 9'b10001010;
				8'b100011: c <= 9'b11110011;
				8'b1110101: c <= 9'b1010001;
				8'b1111101: c <= 9'b100111101;
				8'b101001: c <= 9'b11001101;
				8'b1010010: c <= 9'b11001011;
				8'b1011000: c <= 9'b110001000;
				8'b101110: c <= 9'b110100101;
				8'b1000001: c <= 9'b1101001;
				default: c <= 9'b0;
			endcase
			9'b10111110 : case(di)
				8'b1000011: c <= 9'b101101;
				8'b101000: c <= 9'b11110010;
				8'b111010: c <= 9'b110110010;
				8'b110110: c <= 9'b110100000;
				8'b1100100: c <= 9'b110100111;
				8'b1000000: c <= 9'b110010100;
				8'b1110110: c <= 9'b10001001;
				8'b100101: c <= 9'b1100111;
				8'b101111: c <= 9'b11010;
				8'b100110: c <= 9'b110110110;
				8'b1100011: c <= 9'b111001;
				8'b1001000: c <= 9'b101101001;
				8'b111000: c <= 9'b101110110;
				8'b110001: c <= 9'b100011001;
				8'b1010111: c <= 9'b110011001;
				8'b1001110: c <= 9'b100110100;
				8'b1101010: c <= 9'b110010110;
				8'b1001001: c <= 9'b110010011;
				8'b1100000: c <= 9'b10011001;
				8'b110111: c <= 9'b101011000;
				8'b1011101: c <= 9'b100000111;
				8'b1011011: c <= 9'b111101001;
				8'b111001: c <= 9'b111010100;
				8'b1001010: c <= 9'b111000;
				8'b110011: c <= 9'b110100011;
				8'b1101100: c <= 9'b10010110;
				8'b1110111: c <= 9'b111011010;
				8'b101011: c <= 9'b11001011;
				8'b1101011: c <= 9'b100111100;
				8'b111100: c <= 9'b1000010;
				8'b1000111: c <= 9'b100011100;
				8'b1011111: c <= 9'b101010101;
				8'b1110100: c <= 9'b1110101;
				8'b101101: c <= 9'b1001011;
				8'b1010011: c <= 9'b10101011;
				8'b1100001: c <= 9'b101110110;
				8'b110101: c <= 9'b111101;
				8'b1000100: c <= 9'b11001001;
				8'b1010001: c <= 9'b100;
				8'b1010100: c <= 9'b101001001;
				8'b1100110: c <= 9'b100101;
				8'b101010: c <= 9'b101001110;
				8'b1011110: c <= 9'b11100111;
				8'b1100111: c <= 9'b10010111;
				8'b1011010: c <= 9'b100010;
				8'b1000010: c <= 9'b1100010;
				8'b111101: c <= 9'b11010101;
				8'b110000: c <= 9'b101110001;
				8'b111110: c <= 9'b11000;
				8'b1100010: c <= 9'b10100111;
				8'b1110000: c <= 9'b1000001;
				8'b1101001: c <= 9'b101011011;
				8'b1110011: c <= 9'b111001110;
				8'b1001100: c <= 9'b11011010;
				8'b100001: c <= 9'b11000111;
				8'b1000110: c <= 9'b11010100;
				8'b1110010: c <= 9'b11010011;
				8'b1010000: c <= 9'b1111110;
				8'b1111010: c <= 9'b10001110;
				8'b1010101: c <= 9'b101111001;
				8'b111011: c <= 9'b10000011;
				8'b1001101: c <= 9'b111011001;
				8'b111111: c <= 9'b100000010;
				8'b1101110: c <= 9'b1110000;
				8'b1111011: c <= 9'b11111000;
				8'b1001011: c <= 9'b100101111;
				8'b1101111: c <= 9'b111101000;
				8'b1101000: c <= 9'b11111;
				8'b101100: c <= 9'b111011001;
				8'b100100: c <= 9'b11010011;
				8'b1111000: c <= 9'b100111011;
				8'b1000101: c <= 9'b1011010;
				8'b1011001: c <= 9'b100101001;
				8'b110100: c <= 9'b10000110;
				8'b1111001: c <= 9'b111111110;
				8'b1110001: c <= 9'b101010011;
				8'b1001111: c <= 9'b110011100;
				8'b1100101: c <= 9'b110110110;
				8'b1111110: c <= 9'b10111011;
				8'b1111100: c <= 9'b101100000;
				8'b1010110: c <= 9'b110111111;
				8'b110010: c <= 9'b111011100;
				8'b1101101: c <= 9'b100111010;
				8'b100011: c <= 9'b111000010;
				8'b1110101: c <= 9'b11110011;
				8'b1111101: c <= 9'b10111100;
				8'b101001: c <= 9'b100101;
				8'b1010010: c <= 9'b111100001;
				8'b1011000: c <= 9'b1000101;
				8'b101110: c <= 9'b10010011;
				8'b1000001: c <= 9'b101000101;
				default: c <= 9'b0;
			endcase
			9'b101010101 : case(di)
				8'b1000011: c <= 9'b100001010;
				8'b101000: c <= 9'b110001110;
				8'b111010: c <= 9'b110100001;
				8'b110110: c <= 9'b11111000;
				8'b1100100: c <= 9'b11111101;
				8'b1000000: c <= 9'b10110;
				8'b1110110: c <= 9'b10010011;
				8'b100101: c <= 9'b101000110;
				8'b101111: c <= 9'b111000100;
				8'b100110: c <= 9'b101110010;
				8'b1100011: c <= 9'b100100111;
				8'b1001000: c <= 9'b1000101;
				8'b111000: c <= 9'b110111111;
				8'b110001: c <= 9'b11110011;
				8'b1010111: c <= 9'b110110010;
				8'b1001110: c <= 9'b100011101;
				8'b1101010: c <= 9'b100010000;
				8'b1001001: c <= 9'b101101001;
				8'b1100000: c <= 9'b110011001;
				8'b110111: c <= 9'b11001110;
				8'b1011101: c <= 9'b111001;
				8'b1011011: c <= 9'b100010111;
				8'b111001: c <= 9'b100101011;
				8'b1001010: c <= 9'b11110101;
				8'b110011: c <= 9'b100111100;
				8'b1101100: c <= 9'b11101011;
				8'b1110111: c <= 9'b100111;
				8'b101011: c <= 9'b101110111;
				8'b1101011: c <= 9'b110001110;
				8'b111100: c <= 9'b101110011;
				8'b1000111: c <= 9'b100011111;
				8'b1011111: c <= 9'b110110010;
				8'b1110100: c <= 9'b111000000;
				8'b101101: c <= 9'b101011000;
				8'b1010011: c <= 9'b111110110;
				8'b1100001: c <= 9'b110010;
				8'b110101: c <= 9'b101011010;
				8'b1000100: c <= 9'b10001100;
				8'b1010001: c <= 9'b1011011;
				8'b1010100: c <= 9'b111010110;
				8'b1100110: c <= 9'b1110111;
				8'b101010: c <= 9'b10101011;
				8'b1011110: c <= 9'b111000101;
				8'b1100111: c <= 9'b110010010;
				8'b1011010: c <= 9'b111011101;
				8'b1000010: c <= 9'b101011011;
				8'b111101: c <= 9'b1000110;
				8'b110000: c <= 9'b11010000;
				8'b111110: c <= 9'b10001001;
				8'b1100010: c <= 9'b110001000;
				8'b1110000: c <= 9'b101110001;
				8'b1101001: c <= 9'b10111100;
				8'b1110011: c <= 9'b101001001;
				8'b1001100: c <= 9'b110110010;
				8'b100001: c <= 9'b101100110;
				8'b1000110: c <= 9'b110000000;
				8'b1110010: c <= 9'b100011000;
				8'b1010000: c <= 9'b110101111;
				8'b1111010: c <= 9'b11101011;
				8'b1010101: c <= 9'b11100100;
				8'b111011: c <= 9'b101100001;
				8'b1001101: c <= 9'b101000110;
				8'b111111: c <= 9'b111000111;
				8'b1101110: c <= 9'b1001010;
				8'b1111011: c <= 9'b11100001;
				8'b1001011: c <= 9'b100110111;
				8'b1101111: c <= 9'b111001111;
				8'b1101000: c <= 9'b110101011;
				8'b101100: c <= 9'b1100111;
				8'b100100: c <= 9'b1;
				8'b1111000: c <= 9'b1;
				8'b1000101: c <= 9'b110001110;
				8'b1011001: c <= 9'b1000010;
				8'b110100: c <= 9'b1001111;
				8'b1111001: c <= 9'b1110111;
				8'b1110001: c <= 9'b110110011;
				8'b1001111: c <= 9'b100110100;
				8'b1100101: c <= 9'b101100110;
				8'b1111110: c <= 9'b111011100;
				8'b1111100: c <= 9'b111011001;
				8'b1010110: c <= 9'b1000101;
				8'b110010: c <= 9'b101101001;
				8'b1101101: c <= 9'b1101000;
				8'b100011: c <= 9'b11110101;
				8'b1110101: c <= 9'b101111010;
				8'b1111101: c <= 9'b1010101;
				8'b101001: c <= 9'b11000111;
				8'b1010010: c <= 9'b100010011;
				8'b1011000: c <= 9'b100100011;
				8'b101110: c <= 9'b11100011;
				8'b1000001: c <= 9'b101000001;
				default: c <= 9'b0;
			endcase
			9'b101110100 : case(di)
				8'b1000011: c <= 9'b100001111;
				8'b101000: c <= 9'b101111000;
				8'b111010: c <= 9'b101100101;
				8'b110110: c <= 9'b100110000;
				8'b1100100: c <= 9'b1001110;
				8'b1000000: c <= 9'b111100;
				8'b1110110: c <= 9'b1111101;
				8'b100101: c <= 9'b100010110;
				8'b101111: c <= 9'b100111000;
				8'b100110: c <= 9'b101000;
				8'b1100011: c <= 9'b100100010;
				8'b1001000: c <= 9'b100000001;
				8'b111000: c <= 9'b11001110;
				8'b110001: c <= 9'b110101010;
				8'b1010111: c <= 9'b1111110;
				8'b1001110: c <= 9'b101111001;
				8'b1101010: c <= 9'b111011101;
				8'b1001001: c <= 9'b10100100;
				8'b1100000: c <= 9'b100111010;
				8'b110111: c <= 9'b1110101;
				8'b1011101: c <= 9'b110101100;
				8'b1011011: c <= 9'b101100111;
				8'b111001: c <= 9'b100001011;
				8'b1001010: c <= 9'b101101111;
				8'b110011: c <= 9'b11100100;
				8'b1101100: c <= 9'b100111;
				8'b1110111: c <= 9'b10111000;
				8'b101011: c <= 9'b10101100;
				8'b1101011: c <= 9'b110101101;
				8'b111100: c <= 9'b11100001;
				8'b1000111: c <= 9'b10111111;
				8'b1011111: c <= 9'b11100101;
				8'b1110100: c <= 9'b11110011;
				8'b101101: c <= 9'b11101;
				8'b1010011: c <= 9'b111010010;
				8'b1100001: c <= 9'b111011011;
				8'b110101: c <= 9'b100010011;
				8'b1000100: c <= 9'b1011100;
				8'b1010001: c <= 9'b10011001;
				8'b1010100: c <= 9'b101011001;
				8'b1100110: c <= 9'b10101110;
				8'b101010: c <= 9'b1101110;
				8'b1011110: c <= 9'b110011110;
				8'b1100111: c <= 9'b11100000;
				8'b1011010: c <= 9'b10011010;
				8'b1000010: c <= 9'b110000;
				8'b111101: c <= 9'b100101010;
				8'b110000: c <= 9'b10000011;
				8'b111110: c <= 9'b10111010;
				8'b1100010: c <= 9'b1010000;
				8'b1110000: c <= 9'b110000;
				8'b1101001: c <= 9'b111011110;
				8'b1110011: c <= 9'b110001100;
				8'b1001100: c <= 9'b10011100;
				8'b100001: c <= 9'b111100;
				8'b1000110: c <= 9'b1010010;
				8'b1110010: c <= 9'b1101000;
				8'b1010000: c <= 9'b110001010;
				8'b1111010: c <= 9'b111000010;
				8'b1010101: c <= 9'b100101010;
				8'b111011: c <= 9'b1100011;
				8'b1001101: c <= 9'b1010111;
				8'b111111: c <= 9'b110111111;
				8'b1101110: c <= 9'b111011010;
				8'b1111011: c <= 9'b110000000;
				8'b1001011: c <= 9'b100010010;
				8'b1101111: c <= 9'b111111001;
				8'b1101000: c <= 9'b111001110;
				8'b101100: c <= 9'b100010111;
				8'b100100: c <= 9'b100010011;
				8'b1111000: c <= 9'b10010111;
				8'b1000101: c <= 9'b110100000;
				8'b1011001: c <= 9'b110100110;
				8'b110100: c <= 9'b111100110;
				8'b1111001: c <= 9'b111011100;
				8'b1110001: c <= 9'b110111000;
				8'b1001111: c <= 9'b10000011;
				8'b1100101: c <= 9'b11111;
				8'b1111110: c <= 9'b1100101;
				8'b1111100: c <= 9'b110101101;
				8'b1010110: c <= 9'b100111100;
				8'b110010: c <= 9'b110101111;
				8'b1101101: c <= 9'b1110010;
				8'b100011: c <= 9'b100010010;
				8'b1110101: c <= 9'b11101;
				8'b1111101: c <= 9'b111101110;
				8'b101001: c <= 9'b101001011;
				8'b1010010: c <= 9'b100101111;
				8'b1011000: c <= 9'b101001;
				8'b101110: c <= 9'b111111111;
				8'b1000001: c <= 9'b100110110;
				default: c <= 9'b0;
			endcase
			9'b10100111 : case(di)
				8'b1000011: c <= 9'b110011100;
				8'b101000: c <= 9'b10;
				8'b111010: c <= 9'b101110010;
				8'b110110: c <= 9'b10010011;
				8'b1100100: c <= 9'b111001110;
				8'b1000000: c <= 9'b110100111;
				8'b1110110: c <= 9'b11001001;
				8'b100101: c <= 9'b11010010;
				8'b101111: c <= 9'b11101011;
				8'b100110: c <= 9'b101110011;
				8'b1100011: c <= 9'b10111011;
				8'b1001000: c <= 9'b111011110;
				8'b111000: c <= 9'b110100101;
				8'b110001: c <= 9'b100111101;
				8'b1010111: c <= 9'b111110011;
				8'b1001110: c <= 9'b110011101;
				8'b1101010: c <= 9'b11111001;
				8'b1001001: c <= 9'b10011;
				8'b1100000: c <= 9'b100011010;
				8'b110111: c <= 9'b11110001;
				8'b1011101: c <= 9'b110111100;
				8'b1011011: c <= 9'b10001011;
				8'b111001: c <= 9'b10011001;
				8'b1001010: c <= 9'b101010111;
				8'b110011: c <= 9'b1001010;
				8'b1101100: c <= 9'b100101001;
				8'b1110111: c <= 9'b11;
				8'b101011: c <= 9'b111100111;
				8'b1101011: c <= 9'b10100010;
				8'b111100: c <= 9'b10001011;
				8'b1000111: c <= 9'b110011100;
				8'b1011111: c <= 9'b10011111;
				8'b1110100: c <= 9'b11101100;
				8'b101101: c <= 9'b10100011;
				8'b1010011: c <= 9'b111011;
				8'b1100001: c <= 9'b100111010;
				8'b110101: c <= 9'b100101;
				8'b1000100: c <= 9'b100010000;
				8'b1010001: c <= 9'b111111011;
				8'b1010100: c <= 9'b101011111;
				8'b1100110: c <= 9'b10001101;
				8'b101010: c <= 9'b100000100;
				8'b1011110: c <= 9'b101110001;
				8'b1100111: c <= 9'b10001101;
				8'b1011010: c <= 9'b1101111;
				8'b1000010: c <= 9'b110110000;
				8'b111101: c <= 9'b100111111;
				8'b110000: c <= 9'b10000000;
				8'b111110: c <= 9'b100110110;
				8'b1100010: c <= 9'b100110010;
				8'b1110000: c <= 9'b1001000;
				8'b1101001: c <= 9'b110100010;
				8'b1110011: c <= 9'b10000011;
				8'b1001100: c <= 9'b11001;
				8'b100001: c <= 9'b10101111;
				8'b1000110: c <= 9'b10110011;
				8'b1110010: c <= 9'b111010;
				8'b1010000: c <= 9'b111001111;
				8'b1111010: c <= 9'b11010010;
				8'b1010101: c <= 9'b100101011;
				8'b111011: c <= 9'b1011001;
				8'b1001101: c <= 9'b111100;
				8'b111111: c <= 9'b100001;
				8'b1101110: c <= 9'b110101110;
				8'b1111011: c <= 9'b100111;
				8'b1001011: c <= 9'b111000;
				8'b1101111: c <= 9'b111001001;
				8'b1101000: c <= 9'b1101111;
				8'b101100: c <= 9'b111001011;
				8'b100100: c <= 9'b100100001;
				8'b1111000: c <= 9'b110111111;
				8'b1000101: c <= 9'b110111010;
				8'b1011001: c <= 9'b11011000;
				8'b110100: c <= 9'b10110;
				8'b1111001: c <= 9'b10001010;
				8'b1110001: c <= 9'b110000010;
				8'b1001111: c <= 9'b110110;
				8'b1100101: c <= 9'b11001000;
				8'b1111110: c <= 9'b11111000;
				8'b1111100: c <= 9'b110100111;
				8'b1010110: c <= 9'b10111011;
				8'b110010: c <= 9'b101000001;
				8'b1101101: c <= 9'b1011000;
				8'b100011: c <= 9'b100100010;
				8'b1110101: c <= 9'b10000001;
				8'b1111101: c <= 9'b101101100;
				8'b101001: c <= 9'b111000110;
				8'b1010010: c <= 9'b100;
				8'b1011000: c <= 9'b110010111;
				8'b101110: c <= 9'b1101001;
				8'b1000001: c <= 9'b1001011;
				default: c <= 9'b0;
			endcase
			9'b1011111 : case(di)
				8'b1000011: c <= 9'b1101100;
				8'b101000: c <= 9'b110000110;
				8'b111010: c <= 9'b1000011;
				8'b110110: c <= 9'b1111010;
				8'b1100100: c <= 9'b101011010;
				8'b1000000: c <= 9'b11010100;
				8'b1110110: c <= 9'b100101101;
				8'b100101: c <= 9'b100011100;
				8'b101111: c <= 9'b1110011;
				8'b100110: c <= 9'b100111010;
				8'b1100011: c <= 9'b11100111;
				8'b1001000: c <= 9'b1001110;
				8'b111000: c <= 9'b1000011;
				8'b110001: c <= 9'b110101001;
				8'b1010111: c <= 9'b101111111;
				8'b1001110: c <= 9'b11010100;
				8'b1101010: c <= 9'b1010001;
				8'b1001001: c <= 9'b1000100;
				8'b1100000: c <= 9'b101011010;
				8'b110111: c <= 9'b1000000;
				8'b1011101: c <= 9'b100110000;
				8'b1011011: c <= 9'b100111101;
				8'b111001: c <= 9'b110011011;
				8'b1001010: c <= 9'b101000010;
				8'b110011: c <= 9'b111100000;
				8'b1101100: c <= 9'b10101001;
				8'b1110111: c <= 9'b11110010;
				8'b101011: c <= 9'b111011101;
				8'b1101011: c <= 9'b111001000;
				8'b111100: c <= 9'b101101100;
				8'b1000111: c <= 9'b10100111;
				8'b1011111: c <= 9'b100110100;
				8'b1110100: c <= 9'b1100010;
				8'b101101: c <= 9'b110100;
				8'b1010011: c <= 9'b101110101;
				8'b1100001: c <= 9'b101111000;
				8'b110101: c <= 9'b1011000;
				8'b1000100: c <= 9'b110001;
				8'b1010001: c <= 9'b10011000;
				8'b1010100: c <= 9'b101010100;
				8'b1100110: c <= 9'b110110111;
				8'b101010: c <= 9'b11100100;
				8'b1011110: c <= 9'b101100010;
				8'b1100111: c <= 9'b10111010;
				8'b1011010: c <= 9'b101100110;
				8'b1000010: c <= 9'b10011000;
				8'b111101: c <= 9'b1111;
				8'b110000: c <= 9'b100110;
				8'b111110: c <= 9'b101000110;
				8'b1100010: c <= 9'b101110111;
				8'b1110000: c <= 9'b101010110;
				8'b1101001: c <= 9'b10011000;
				8'b1110011: c <= 9'b1000001;
				8'b1001100: c <= 9'b111101111;
				8'b100001: c <= 9'b101000001;
				8'b1000110: c <= 9'b100110110;
				8'b1110010: c <= 9'b10010000;
				8'b1010000: c <= 9'b1100000;
				8'b1111010: c <= 9'b100111100;
				8'b1010101: c <= 9'b110010101;
				8'b111011: c <= 9'b10000;
				8'b1001101: c <= 9'b111010001;
				8'b111111: c <= 9'b11011101;
				8'b1101110: c <= 9'b110111011;
				8'b1111011: c <= 9'b101000011;
				8'b1001011: c <= 9'b100101001;
				8'b1101111: c <= 9'b100001011;
				8'b1101000: c <= 9'b100000100;
				8'b101100: c <= 9'b100001010;
				8'b100100: c <= 9'b11001;
				8'b1111000: c <= 9'b1001;
				8'b1000101: c <= 9'b10000110;
				8'b1011001: c <= 9'b110011100;
				8'b110100: c <= 9'b100011010;
				8'b1111001: c <= 9'b10001110;
				8'b1110001: c <= 9'b110010001;
				8'b1001111: c <= 9'b10011100;
				8'b1100101: c <= 9'b111000101;
				8'b1111110: c <= 9'b101110101;
				8'b1111100: c <= 9'b10110011;
				8'b1010110: c <= 9'b1011011;
				8'b110010: c <= 9'b110101011;
				8'b1101101: c <= 9'b100000001;
				8'b100011: c <= 9'b101110110;
				8'b1110101: c <= 9'b110011111;
				8'b1111101: c <= 9'b1100101;
				8'b101001: c <= 9'b110000000;
				8'b1010010: c <= 9'b101100100;
				8'b1011000: c <= 9'b11000111;
				8'b101110: c <= 9'b1001010;
				8'b1000001: c <= 9'b110100100;
				default: c <= 9'b0;
			endcase
			9'b101100001 : case(di)
				8'b1000011: c <= 9'b100100101;
				8'b101000: c <= 9'b101100;
				8'b111010: c <= 9'b1111;
				8'b110110: c <= 9'b100101101;
				8'b1100100: c <= 9'b1000001;
				8'b1000000: c <= 9'b100101111;
				8'b1110110: c <= 9'b100101011;
				8'b100101: c <= 9'b110100110;
				8'b101111: c <= 9'b11100111;
				8'b100110: c <= 9'b10111011;
				8'b1100011: c <= 9'b101000001;
				8'b1001000: c <= 9'b111001001;
				8'b111000: c <= 9'b11010;
				8'b110001: c <= 9'b10001110;
				8'b1010111: c <= 9'b100110000;
				8'b1001110: c <= 9'b100010101;
				8'b1101010: c <= 9'b101101000;
				8'b1001001: c <= 9'b101001111;
				8'b1100000: c <= 9'b111100101;
				8'b110111: c <= 9'b100;
				8'b1011101: c <= 9'b10101001;
				8'b1011011: c <= 9'b10000011;
				8'b111001: c <= 9'b100111010;
				8'b1001010: c <= 9'b110111100;
				8'b110011: c <= 9'b10110100;
				8'b1101100: c <= 9'b10001000;
				8'b1110111: c <= 9'b10111100;
				8'b101011: c <= 9'b11111000;
				8'b1101011: c <= 9'b1100101;
				8'b111100: c <= 9'b100100;
				8'b1000111: c <= 9'b110100001;
				8'b1011111: c <= 9'b101100010;
				8'b1110100: c <= 9'b10111;
				8'b101101: c <= 9'b101110110;
				8'b1010011: c <= 9'b101000100;
				8'b1100001: c <= 9'b101111110;
				8'b110101: c <= 9'b110110110;
				8'b1000100: c <= 9'b10101111;
				8'b1010001: c <= 9'b111000111;
				8'b1010100: c <= 9'b10011001;
				8'b1100110: c <= 9'b111001110;
				8'b101010: c <= 9'b10001000;
				8'b1011110: c <= 9'b1010111;
				8'b1100111: c <= 9'b111010;
				8'b1011010: c <= 9'b110001011;
				8'b1000010: c <= 9'b110001100;
				8'b111101: c <= 9'b110111111;
				8'b110000: c <= 9'b101;
				8'b111110: c <= 9'b100001111;
				8'b1100010: c <= 9'b101000001;
				8'b1110000: c <= 9'b111010010;
				8'b1101001: c <= 9'b101110;
				8'b1110011: c <= 9'b101000010;
				8'b1001100: c <= 9'b10000110;
				8'b100001: c <= 9'b10010001;
				8'b1000110: c <= 9'b11010;
				8'b1110010: c <= 9'b10110101;
				8'b1010000: c <= 9'b100101;
				8'b1111010: c <= 9'b11000010;
				8'b1010101: c <= 9'b101010111;
				8'b111011: c <= 9'b101111111;
				8'b1001101: c <= 9'b100101110;
				8'b111111: c <= 9'b11011010;
				8'b1101110: c <= 9'b101001011;
				8'b1111011: c <= 9'b110010101;
				8'b1001011: c <= 9'b100001100;
				8'b1101111: c <= 9'b1000000;
				8'b1101000: c <= 9'b11111001;
				8'b101100: c <= 9'b100011011;
				8'b100100: c <= 9'b10010101;
				8'b1111000: c <= 9'b110100010;
				8'b1000101: c <= 9'b11000010;
				8'b1011001: c <= 9'b11000001;
				8'b110100: c <= 9'b10010101;
				8'b1111001: c <= 9'b11001000;
				8'b1110001: c <= 9'b1111001;
				8'b1001111: c <= 9'b10101101;
				8'b1100101: c <= 9'b1110010;
				8'b1111110: c <= 9'b10111100;
				8'b1111100: c <= 9'b10100111;
				8'b1010110: c <= 9'b110101110;
				8'b110010: c <= 9'b11100101;
				8'b1101101: c <= 9'b110001101;
				8'b100011: c <= 9'b101100101;
				8'b1110101: c <= 9'b100110;
				8'b1111101: c <= 9'b100110111;
				8'b101001: c <= 9'b111100001;
				8'b1010010: c <= 9'b100101110;
				8'b1011000: c <= 9'b10111000;
				8'b101110: c <= 9'b111010110;
				8'b1000001: c <= 9'b1010111;
				default: c <= 9'b0;
			endcase
			9'b11010 : case(di)
				8'b1000011: c <= 9'b10010111;
				8'b101000: c <= 9'b100111100;
				8'b111010: c <= 9'b11101000;
				8'b110110: c <= 9'b101100;
				8'b1100100: c <= 9'b100011100;
				8'b1000000: c <= 9'b100100001;
				8'b1110110: c <= 9'b100100010;
				8'b100101: c <= 9'b101010100;
				8'b101111: c <= 9'b10010101;
				8'b100110: c <= 9'b100110000;
				8'b1100011: c <= 9'b101110010;
				8'b1001000: c <= 9'b110000010;
				8'b111000: c <= 9'b1011100;
				8'b110001: c <= 9'b1111011;
				8'b1010111: c <= 9'b111010110;
				8'b1001110: c <= 9'b11001110;
				8'b1101010: c <= 9'b110110100;
				8'b1001001: c <= 9'b101011001;
				8'b1100000: c <= 9'b11001100;
				8'b110111: c <= 9'b110011011;
				8'b1011101: c <= 9'b11010100;
				8'b1011011: c <= 9'b100010110;
				8'b111001: c <= 9'b1100100;
				8'b1001010: c <= 9'b11000111;
				8'b110011: c <= 9'b110111;
				8'b1101100: c <= 9'b1100101;
				8'b1110111: c <= 9'b10010001;
				8'b101011: c <= 9'b111001110;
				8'b1101011: c <= 9'b110011001;
				8'b111100: c <= 9'b100101111;
				8'b1000111: c <= 9'b11011011;
				8'b1011111: c <= 9'b101010110;
				8'b1110100: c <= 9'b111000101;
				8'b101101: c <= 9'b10101011;
				8'b1010011: c <= 9'b10110;
				8'b1100001: c <= 9'b1001100;
				8'b110101: c <= 9'b111011010;
				8'b1000100: c <= 9'b111010010;
				8'b1010001: c <= 9'b11010100;
				8'b1010100: c <= 9'b101001011;
				8'b1100110: c <= 9'b10000110;
				8'b101010: c <= 9'b10100000;
				8'b1011110: c <= 9'b10011101;
				8'b1100111: c <= 9'b101101001;
				8'b1011010: c <= 9'b101000;
				8'b1000010: c <= 9'b11011010;
				8'b111101: c <= 9'b101010101;
				8'b110000: c <= 9'b101001000;
				8'b111110: c <= 9'b10;
				8'b1100010: c <= 9'b111000000;
				8'b1110000: c <= 9'b1001001;
				8'b1101001: c <= 9'b111011001;
				8'b1110011: c <= 9'b100111;
				8'b1001100: c <= 9'b111001001;
				8'b100001: c <= 9'b10100000;
				8'b1000110: c <= 9'b10010000;
				8'b1110010: c <= 9'b110100001;
				8'b1010000: c <= 9'b111011;
				8'b1111010: c <= 9'b11100101;
				8'b1010101: c <= 9'b10001001;
				8'b111011: c <= 9'b111010111;
				8'b1001101: c <= 9'b10100101;
				8'b111111: c <= 9'b100010101;
				8'b1101110: c <= 9'b101101;
				8'b1111011: c <= 9'b101001110;
				8'b1001011: c <= 9'b1000011;
				8'b1101111: c <= 9'b100101001;
				8'b1101000: c <= 9'b101100100;
				8'b101100: c <= 9'b11101111;
				8'b100100: c <= 9'b1000001;
				8'b1111000: c <= 9'b10000011;
				8'b1000101: c <= 9'b10101101;
				8'b1011001: c <= 9'b10000;
				8'b110100: c <= 9'b11011110;
				8'b1111001: c <= 9'b101001010;
				8'b1110001: c <= 9'b111011101;
				8'b1001111: c <= 9'b1010000;
				8'b1100101: c <= 9'b101000101;
				8'b1111110: c <= 9'b10101111;
				8'b1111100: c <= 9'b100011011;
				8'b1010110: c <= 9'b1001110;
				8'b110010: c <= 9'b100111;
				8'b1101101: c <= 9'b111001010;
				8'b100011: c <= 9'b10100111;
				8'b1110101: c <= 9'b1101;
				8'b1111101: c <= 9'b110100000;
				8'b101001: c <= 9'b110111001;
				8'b1010010: c <= 9'b111000000;
				8'b1011000: c <= 9'b101101101;
				8'b101110: c <= 9'b111011;
				8'b1000001: c <= 9'b100010010;
				default: c <= 9'b0;
			endcase
			9'b110001111 : case(di)
				8'b1000011: c <= 9'b110011111;
				8'b101000: c <= 9'b100101;
				8'b111010: c <= 9'b111000000;
				8'b110110: c <= 9'b111100101;
				8'b1100100: c <= 9'b101100100;
				8'b1000000: c <= 9'b10010111;
				8'b1110110: c <= 9'b1111;
				8'b100101: c <= 9'b110001000;
				8'b101111: c <= 9'b101100101;
				8'b100110: c <= 9'b100011101;
				8'b1100011: c <= 9'b111111000;
				8'b1001000: c <= 9'b101111000;
				8'b111000: c <= 9'b100010;
				8'b110001: c <= 9'b10001010;
				8'b1010111: c <= 9'b11111000;
				8'b1001110: c <= 9'b111;
				8'b1101010: c <= 9'b101101100;
				8'b1001001: c <= 9'b110110010;
				8'b1100000: c <= 9'b100000010;
				8'b110111: c <= 9'b111000;
				8'b1011101: c <= 9'b1110100;
				8'b1011011: c <= 9'b111011110;
				8'b111001: c <= 9'b10011101;
				8'b1001010: c <= 9'b110000;
				8'b110011: c <= 9'b1111111;
				8'b1101100: c <= 9'b10000101;
				8'b1110111: c <= 9'b111001;
				8'b101011: c <= 9'b110101010;
				8'b1101011: c <= 9'b101011111;
				8'b111100: c <= 9'b110011101;
				8'b1000111: c <= 9'b1110001;
				8'b1011111: c <= 9'b110000101;
				8'b1110100: c <= 9'b111000100;
				8'b101101: c <= 9'b11010101;
				8'b1010011: c <= 9'b111001100;
				8'b1100001: c <= 9'b110001011;
				8'b110101: c <= 9'b111100101;
				8'b1000100: c <= 9'b1001001;
				8'b1010001: c <= 9'b111110101;
				8'b1010100: c <= 9'b10100010;
				8'b1100110: c <= 9'b11010101;
				8'b101010: c <= 9'b101101100;
				8'b1011110: c <= 9'b100100001;
				8'b1100111: c <= 9'b101010001;
				8'b1011010: c <= 9'b110101;
				8'b1000010: c <= 9'b101101001;
				8'b111101: c <= 9'b111010010;
				8'b110000: c <= 9'b110100010;
				8'b111110: c <= 9'b110001110;
				8'b1100010: c <= 9'b11111110;
				8'b1110000: c <= 9'b11001011;
				8'b1101001: c <= 9'b11010101;
				8'b1110011: c <= 9'b110001;
				8'b1001100: c <= 9'b1110011;
				8'b100001: c <= 9'b110101110;
				8'b1000110: c <= 9'b100010011;
				8'b1110010: c <= 9'b111010010;
				8'b1010000: c <= 9'b110101100;
				8'b1111010: c <= 9'b100011111;
				8'b1010101: c <= 9'b11101000;
				8'b111011: c <= 9'b110001;
				8'b1001101: c <= 9'b110100111;
				8'b111111: c <= 9'b1100100;
				8'b1101110: c <= 9'b110010010;
				8'b1111011: c <= 9'b1001;
				8'b1001011: c <= 9'b100101000;
				8'b1101111: c <= 9'b100010001;
				8'b1101000: c <= 9'b101010011;
				8'b101100: c <= 9'b100110100;
				8'b100100: c <= 9'b11110011;
				8'b1111000: c <= 9'b110110010;
				8'b1000101: c <= 9'b100011100;
				8'b1011001: c <= 9'b11000001;
				8'b110100: c <= 9'b100100000;
				8'b1111001: c <= 9'b111111010;
				8'b1110001: c <= 9'b110000000;
				8'b1001111: c <= 9'b101011110;
				8'b1100101: c <= 9'b11101101;
				8'b1111110: c <= 9'b1100101;
				8'b1111100: c <= 9'b1000010;
				8'b1010110: c <= 9'b111110001;
				8'b110010: c <= 9'b11011101;
				8'b1101101: c <= 9'b110000;
				8'b100011: c <= 9'b101000110;
				8'b1110101: c <= 9'b110010011;
				8'b1111101: c <= 9'b1011100;
				8'b101001: c <= 9'b100010000;
				8'b1010010: c <= 9'b1101001;
				8'b1011000: c <= 9'b111111110;
				8'b101110: c <= 9'b111001001;
				8'b1000001: c <= 9'b111111111;
				default: c <= 9'b0;
			endcase
			9'b11101000 : case(di)
				8'b1000011: c <= 9'b11100110;
				8'b101000: c <= 9'b100011000;
				8'b111010: c <= 9'b1011001;
				8'b110110: c <= 9'b110110100;
				8'b1100100: c <= 9'b110111001;
				8'b1000000: c <= 9'b101011001;
				8'b1110110: c <= 9'b110110111;
				8'b100101: c <= 9'b100100001;
				8'b101111: c <= 9'b11000111;
				8'b100110: c <= 9'b100101110;
				8'b1100011: c <= 9'b10010110;
				8'b1001000: c <= 9'b100101001;
				8'b111000: c <= 9'b110111111;
				8'b110001: c <= 9'b11010111;
				8'b1010111: c <= 9'b111010111;
				8'b1001110: c <= 9'b101111000;
				8'b1101010: c <= 9'b11101000;
				8'b1001001: c <= 9'b11101111;
				8'b1100000: c <= 9'b110010100;
				8'b110111: c <= 9'b100111000;
				8'b1011101: c <= 9'b100010011;
				8'b1011011: c <= 9'b100000111;
				8'b111001: c <= 9'b1010011;
				8'b1001010: c <= 9'b1010001;
				8'b110011: c <= 9'b111010001;
				8'b1101100: c <= 9'b100111;
				8'b1110111: c <= 9'b1110001;
				8'b101011: c <= 9'b110100011;
				8'b1101011: c <= 9'b11110001;
				8'b111100: c <= 9'b110001010;
				8'b1000111: c <= 9'b110011111;
				8'b1011111: c <= 9'b111101001;
				8'b1110100: c <= 9'b101101110;
				8'b101101: c <= 9'b10001110;
				8'b1010011: c <= 9'b1000001;
				8'b1100001: c <= 9'b10110100;
				8'b110101: c <= 9'b11001;
				8'b1000100: c <= 9'b101011101;
				8'b1010001: c <= 9'b101110001;
				8'b1010100: c <= 9'b11110000;
				8'b1100110: c <= 9'b10001100;
				8'b101010: c <= 9'b100100110;
				8'b1011110: c <= 9'b100110;
				8'b1100111: c <= 9'b110101111;
				8'b1011010: c <= 9'b110100;
				8'b1000010: c <= 9'b11011;
				8'b111101: c <= 9'b10000001;
				8'b110000: c <= 9'b101000010;
				8'b111110: c <= 9'b11110001;
				8'b1100010: c <= 9'b10110;
				8'b1110000: c <= 9'b110001000;
				8'b1101001: c <= 9'b101101001;
				8'b1110011: c <= 9'b1111001;
				8'b1001100: c <= 9'b10100;
				8'b100001: c <= 9'b110001011;
				8'b1000110: c <= 9'b101001001;
				8'b1110010: c <= 9'b100110110;
				8'b1010000: c <= 9'b11000001;
				8'b1111010: c <= 9'b110100100;
				8'b1010101: c <= 9'b11011110;
				8'b111011: c <= 9'b11110110;
				8'b1001101: c <= 9'b111010100;
				8'b111111: c <= 9'b11010000;
				8'b1101110: c <= 9'b11010111;
				8'b1111011: c <= 9'b11011010;
				8'b1001011: c <= 9'b1000101;
				8'b1101111: c <= 9'b111100100;
				8'b1101000: c <= 9'b110010111;
				8'b101100: c <= 9'b10001001;
				8'b100100: c <= 9'b100111011;
				8'b1111000: c <= 9'b1100000;
				8'b1000101: c <= 9'b110001001;
				8'b1011001: c <= 9'b10011100;
				8'b110100: c <= 9'b1001011;
				8'b1111001: c <= 9'b110010100;
				8'b1110001: c <= 9'b11111;
				8'b1001111: c <= 9'b11011010;
				8'b1100101: c <= 9'b110000011;
				8'b1111110: c <= 9'b10000001;
				8'b1111100: c <= 9'b111111000;
				8'b1010110: c <= 9'b111010;
				8'b110010: c <= 9'b111110101;
				8'b1101101: c <= 9'b111110101;
				8'b100011: c <= 9'b111100;
				8'b1110101: c <= 9'b110101001;
				8'b1111101: c <= 9'b1101000;
				8'b101001: c <= 9'b110101110;
				8'b1010010: c <= 9'b100110100;
				8'b1011000: c <= 9'b1011111;
				8'b101110: c <= 9'b11001011;
				8'b1000001: c <= 9'b101110101;
				default: c <= 9'b0;
			endcase
			9'b100011001 : case(di)
				8'b1000011: c <= 9'b11110101;
				8'b101000: c <= 9'b10110;
				8'b111010: c <= 9'b110011010;
				8'b110110: c <= 9'b110001110;
				8'b1100100: c <= 9'b101101011;
				8'b1000000: c <= 9'b110111;
				8'b1110110: c <= 9'b110110010;
				8'b100101: c <= 9'b110001;
				8'b101111: c <= 9'b110111111;
				8'b100110: c <= 9'b101011000;
				8'b1100011: c <= 9'b10101101;
				8'b1001000: c <= 9'b11100110;
				8'b111000: c <= 9'b111111101;
				8'b110001: c <= 9'b100011011;
				8'b1010111: c <= 9'b100001011;
				8'b1001110: c <= 9'b111010000;
				8'b1101010: c <= 9'b101101101;
				8'b1001001: c <= 9'b11111100;
				8'b1100000: c <= 9'b11001011;
				8'b110111: c <= 9'b101000011;
				8'b1011101: c <= 9'b101010011;
				8'b1011011: c <= 9'b1100001;
				8'b111001: c <= 9'b100011000;
				8'b1001010: c <= 9'b11001110;
				8'b110011: c <= 9'b10000101;
				8'b1101100: c <= 9'b110011000;
				8'b1110111: c <= 9'b1000001;
				8'b101011: c <= 9'b11001001;
				8'b1101011: c <= 9'b110010100;
				8'b111100: c <= 9'b101011011;
				8'b1000111: c <= 9'b100011001;
				8'b1011111: c <= 9'b11110010;
				8'b1110100: c <= 9'b100100101;
				8'b101101: c <= 9'b100011;
				8'b1010011: c <= 9'b101010011;
				8'b1100001: c <= 9'b11011011;
				8'b110101: c <= 9'b110110;
				8'b1000100: c <= 9'b1;
				8'b1010001: c <= 9'b111110001;
				8'b1010100: c <= 9'b110110010;
				8'b1100110: c <= 9'b100111111;
				8'b101010: c <= 9'b100000010;
				8'b1011110: c <= 9'b11001;
				8'b1100111: c <= 9'b111111000;
				8'b1011010: c <= 9'b100011010;
				8'b1000010: c <= 9'b110100111;
				8'b111101: c <= 9'b10100;
				8'b110000: c <= 9'b10100000;
				8'b111110: c <= 9'b111110110;
				8'b1100010: c <= 9'b101101101;
				8'b1110000: c <= 9'b1000101;
				8'b1101001: c <= 9'b101011;
				8'b1110011: c <= 9'b10000;
				8'b1001100: c <= 9'b100110101;
				8'b100001: c <= 9'b1001110;
				8'b1000110: c <= 9'b110110111;
				8'b1110010: c <= 9'b100001111;
				8'b1010000: c <= 9'b110100100;
				8'b1111010: c <= 9'b110100;
				8'b1010101: c <= 9'b11010101;
				8'b111011: c <= 9'b11001000;
				8'b1001101: c <= 9'b100001110;
				8'b111111: c <= 9'b111111101;
				8'b1101110: c <= 9'b110000010;
				8'b1111011: c <= 9'b10011101;
				8'b1001011: c <= 9'b100000101;
				8'b1101111: c <= 9'b100111;
				8'b1101000: c <= 9'b11111;
				8'b101100: c <= 9'b1001001;
				8'b100100: c <= 9'b11110111;
				8'b1111000: c <= 9'b1;
				8'b1000101: c <= 9'b111000011;
				8'b1011001: c <= 9'b10110100;
				8'b110100: c <= 9'b10000;
				8'b1111001: c <= 9'b11110;
				8'b1110001: c <= 9'b10001000;
				8'b1001111: c <= 9'b111101100;
				8'b1100101: c <= 9'b101000111;
				8'b1111110: c <= 9'b10010100;
				8'b1111100: c <= 9'b1101111;
				8'b1010110: c <= 9'b1101000;
				8'b110010: c <= 9'b101011111;
				8'b1101101: c <= 9'b10001111;
				8'b100011: c <= 9'b111011110;
				8'b1110101: c <= 9'b110101;
				8'b1111101: c <= 9'b110111;
				8'b101001: c <= 9'b100101010;
				8'b1010010: c <= 9'b11011000;
				8'b1011000: c <= 9'b101101011;
				8'b101110: c <= 9'b101001010;
				8'b1000001: c <= 9'b111011111;
				default: c <= 9'b0;
			endcase
			9'b101010010 : case(di)
				8'b1000011: c <= 9'b10100100;
				8'b101000: c <= 9'b101101111;
				8'b111010: c <= 9'b11000111;
				8'b110110: c <= 9'b100111;
				8'b1100100: c <= 9'b10010;
				8'b1000000: c <= 9'b110000110;
				8'b1110110: c <= 9'b110101101;
				8'b100101: c <= 9'b100110100;
				8'b101111: c <= 9'b100101;
				8'b100110: c <= 9'b111000101;
				8'b1100011: c <= 9'b110000111;
				8'b1001000: c <= 9'b1100110;
				8'b111000: c <= 9'b111111110;
				8'b110001: c <= 9'b101111110;
				8'b1010111: c <= 9'b11001;
				8'b1001110: c <= 9'b110110011;
				8'b1101010: c <= 9'b11101000;
				8'b1001001: c <= 9'b11100111;
				8'b1100000: c <= 9'b10110;
				8'b110111: c <= 9'b111111000;
				8'b1011101: c <= 9'b110001010;
				8'b1011011: c <= 9'b101111010;
				8'b111001: c <= 9'b110101010;
				8'b1001010: c <= 9'b101101010;
				8'b110011: c <= 9'b1000100;
				8'b1101100: c <= 9'b10011001;
				8'b1110111: c <= 9'b1001010;
				8'b101011: c <= 9'b1110010;
				8'b1101011: c <= 9'b11000111;
				8'b111100: c <= 9'b11101111;
				8'b1000111: c <= 9'b1101;
				8'b1011111: c <= 9'b100000101;
				8'b1110100: c <= 9'b100110;
				8'b101101: c <= 9'b110111011;
				8'b1010011: c <= 9'b101100011;
				8'b1100001: c <= 9'b110111000;
				8'b110101: c <= 9'b10100100;
				8'b1000100: c <= 9'b101000100;
				8'b1010001: c <= 9'b101000100;
				8'b1010100: c <= 9'b11101011;
				8'b1100110: c <= 9'b111100010;
				8'b101010: c <= 9'b100000110;
				8'b1011110: c <= 9'b100110010;
				8'b1100111: c <= 9'b1110011;
				8'b1011010: c <= 9'b101101101;
				8'b1000010: c <= 9'b100101011;
				8'b111101: c <= 9'b111100011;
				8'b110000: c <= 9'b10000000;
				8'b111110: c <= 9'b10110111;
				8'b1100010: c <= 9'b100101100;
				8'b1110000: c <= 9'b111000010;
				8'b1101001: c <= 9'b11101;
				8'b1110011: c <= 9'b111000011;
				8'b1001100: c <= 9'b101101011;
				8'b100001: c <= 9'b11010100;
				8'b1000110: c <= 9'b100111011;
				8'b1110010: c <= 9'b101011110;
				8'b1010000: c <= 9'b1000111;
				8'b1111010: c <= 9'b110001000;
				8'b1010101: c <= 9'b11011110;
				8'b111011: c <= 9'b1110100;
				8'b1001101: c <= 9'b100011011;
				8'b111111: c <= 9'b110111110;
				8'b1101110: c <= 9'b111100000;
				8'b1111011: c <= 9'b100010110;
				8'b1001011: c <= 9'b10001000;
				8'b1101111: c <= 9'b110010100;
				8'b1101000: c <= 9'b100111111;
				8'b101100: c <= 9'b101000001;
				8'b100100: c <= 9'b111000010;
				8'b1111000: c <= 9'b100010111;
				8'b1000101: c <= 9'b1110000;
				8'b1011001: c <= 9'b11011000;
				8'b110100: c <= 9'b1111010;
				8'b1111001: c <= 9'b100011;
				8'b1110001: c <= 9'b100010110;
				8'b1001111: c <= 9'b111101000;
				8'b1100101: c <= 9'b10101000;
				8'b1111110: c <= 9'b1001;
				8'b1111100: c <= 9'b110100;
				8'b1010110: c <= 9'b10011111;
				8'b110010: c <= 9'b10001101;
				8'b1101101: c <= 9'b110101101;
				8'b100011: c <= 9'b110001110;
				8'b1110101: c <= 9'b10100100;
				8'b1111101: c <= 9'b100010011;
				8'b101001: c <= 9'b11000100;
				8'b1010010: c <= 9'b100011010;
				8'b1011000: c <= 9'b100110101;
				8'b101110: c <= 9'b110110110;
				8'b1000001: c <= 9'b100100101;
				default: c <= 9'b0;
			endcase
			9'b111011111 : case(di)
				8'b1000011: c <= 9'b1010000;
				8'b101000: c <= 9'b11010100;
				8'b111010: c <= 9'b100101000;
				8'b110110: c <= 9'b101010001;
				8'b1100100: c <= 9'b10110011;
				8'b1000000: c <= 9'b101100011;
				8'b1110110: c <= 9'b100001011;
				8'b100101: c <= 9'b101110111;
				8'b101111: c <= 9'b101001110;
				8'b100110: c <= 9'b1100011;
				8'b1100011: c <= 9'b110101001;
				8'b1001000: c <= 9'b110011111;
				8'b111000: c <= 9'b100010101;
				8'b110001: c <= 9'b101010110;
				8'b1010111: c <= 9'b11001110;
				8'b1001110: c <= 9'b111000101;
				8'b1101010: c <= 9'b101101001;
				8'b1001001: c <= 9'b11001;
				8'b1100000: c <= 9'b11000110;
				8'b110111: c <= 9'b10000011;
				8'b1011101: c <= 9'b101001111;
				8'b1011011: c <= 9'b1001001;
				8'b111001: c <= 9'b111100;
				8'b1001010: c <= 9'b1101110;
				8'b110011: c <= 9'b100011111;
				8'b1101100: c <= 9'b100011100;
				8'b1110111: c <= 9'b1110100;
				8'b101011: c <= 9'b111000110;
				8'b1101011: c <= 9'b11110;
				8'b111100: c <= 9'b111001111;
				8'b1000111: c <= 9'b1000000;
				8'b1011111: c <= 9'b110011101;
				8'b1110100: c <= 9'b111100011;
				8'b101101: c <= 9'b111011;
				8'b1010011: c <= 9'b100101010;
				8'b1100001: c <= 9'b101000001;
				8'b110101: c <= 9'b11001011;
				8'b1000100: c <= 9'b1011100;
				8'b1010001: c <= 9'b11010111;
				8'b1010100: c <= 9'b1000011;
				8'b1100110: c <= 9'b1110111;
				8'b101010: c <= 9'b10111101;
				8'b1011110: c <= 9'b111101001;
				8'b1100111: c <= 9'b111010110;
				8'b1011010: c <= 9'b100111;
				8'b1000010: c <= 9'b11000;
				8'b111101: c <= 9'b111011111;
				8'b110000: c <= 9'b110011000;
				8'b111110: c <= 9'b111010010;
				8'b1100010: c <= 9'b111001011;
				8'b1110000: c <= 9'b10111101;
				8'b1101001: c <= 9'b11100111;
				8'b1110011: c <= 9'b11001101;
				8'b1001100: c <= 9'b1101101;
				8'b100001: c <= 9'b100010;
				8'b1000110: c <= 9'b110110000;
				8'b1110010: c <= 9'b10101001;
				8'b1010000: c <= 9'b11110000;
				8'b1111010: c <= 9'b111011001;
				8'b1010101: c <= 9'b110010100;
				8'b111011: c <= 9'b11010111;
				8'b1001101: c <= 9'b1100;
				8'b111111: c <= 9'b11110100;
				8'b1101110: c <= 9'b100100000;
				8'b1111011: c <= 9'b110010101;
				8'b1001011: c <= 9'b10111011;
				8'b1101111: c <= 9'b10111100;
				8'b1101000: c <= 9'b100100111;
				8'b101100: c <= 9'b10110100;
				8'b100100: c <= 9'b110101001;
				8'b1111000: c <= 9'b11011;
				8'b1000101: c <= 9'b11111010;
				8'b1011001: c <= 9'b100010011;
				8'b110100: c <= 9'b100001001;
				8'b1111001: c <= 9'b101001;
				8'b1110001: c <= 9'b10101000;
				8'b1001111: c <= 9'b11100111;
				8'b1100101: c <= 9'b1011000;
				8'b1111110: c <= 9'b11110010;
				8'b1111100: c <= 9'b11110001;
				8'b1010110: c <= 9'b11010001;
				8'b110010: c <= 9'b110101010;
				8'b1101101: c <= 9'b1111111;
				8'b100011: c <= 9'b110011100;
				8'b1110101: c <= 9'b10010110;
				8'b1111101: c <= 9'b1010110;
				8'b101001: c <= 9'b11010001;
				8'b1010010: c <= 9'b100000110;
				8'b1011000: c <= 9'b110010001;
				8'b101110: c <= 9'b10010110;
				8'b1000001: c <= 9'b10011000;
				default: c <= 9'b0;
			endcase
			9'b11011000 : case(di)
				8'b1000011: c <= 9'b110111;
				8'b101000: c <= 9'b10001011;
				8'b111010: c <= 9'b1000110;
				8'b110110: c <= 9'b11001011;
				8'b1100100: c <= 9'b111000101;
				8'b1000000: c <= 9'b111001001;
				8'b1110110: c <= 9'b11001011;
				8'b100101: c <= 9'b11000110;
				8'b101111: c <= 9'b101110011;
				8'b100110: c <= 9'b10001110;
				8'b1100011: c <= 9'b11101011;
				8'b1001000: c <= 9'b111111011;
				8'b111000: c <= 9'b111000000;
				8'b110001: c <= 9'b10000110;
				8'b1010111: c <= 9'b111101;
				8'b1001110: c <= 9'b111111110;
				8'b1101010: c <= 9'b111100101;
				8'b1001001: c <= 9'b101000111;
				8'b1100000: c <= 9'b11001100;
				8'b110111: c <= 9'b111000011;
				8'b1011101: c <= 9'b101010111;
				8'b1011011: c <= 9'b10001111;
				8'b111001: c <= 9'b100011010;
				8'b1001010: c <= 9'b10001011;
				8'b110011: c <= 9'b101100;
				8'b1101100: c <= 9'b111111;
				8'b1110111: c <= 9'b110001110;
				8'b101011: c <= 9'b11110000;
				8'b1101011: c <= 9'b1101100;
				8'b111100: c <= 9'b101011101;
				8'b1000111: c <= 9'b10010110;
				8'b1011111: c <= 9'b111011;
				8'b1110100: c <= 9'b10101000;
				8'b101101: c <= 9'b11110000;
				8'b1010011: c <= 9'b101000101;
				8'b1100001: c <= 9'b11001011;
				8'b110101: c <= 9'b100101011;
				8'b1000100: c <= 9'b110100110;
				8'b1010001: c <= 9'b100111101;
				8'b1010100: c <= 9'b10111001;
				8'b1100110: c <= 9'b111001000;
				8'b101010: c <= 9'b100100010;
				8'b1011110: c <= 9'b111100;
				8'b1100111: c <= 9'b1100011;
				8'b1011010: c <= 9'b11000011;
				8'b1000010: c <= 9'b1000010;
				8'b111101: c <= 9'b101111001;
				8'b110000: c <= 9'b11011101;
				8'b111110: c <= 9'b1110010;
				8'b1100010: c <= 9'b10001101;
				8'b1110000: c <= 9'b111;
				8'b1101001: c <= 9'b11101011;
				8'b1110011: c <= 9'b1010010;
				8'b1001100: c <= 9'b11000100;
				8'b100001: c <= 9'b1010001;
				8'b1000110: c <= 9'b1000101;
				8'b1110010: c <= 9'b10110101;
				8'b1010000: c <= 9'b1111;
				8'b1111010: c <= 9'b110100101;
				8'b1010101: c <= 9'b111001111;
				8'b111011: c <= 9'b101010110;
				8'b1001101: c <= 9'b100111;
				8'b111111: c <= 9'b110001111;
				8'b1101110: c <= 9'b111101110;
				8'b1111011: c <= 9'b101101101;
				8'b1001011: c <= 9'b101100111;
				8'b1101111: c <= 9'b110110011;
				8'b1101000: c <= 9'b11110110;
				8'b101100: c <= 9'b110011100;
				8'b100100: c <= 9'b110101111;
				8'b1111000: c <= 9'b111000;
				8'b1000101: c <= 9'b111001100;
				8'b1011001: c <= 9'b101101011;
				8'b110100: c <= 9'b101000110;
				8'b1111001: c <= 9'b1110011;
				8'b1110001: c <= 9'b100001110;
				8'b1001111: c <= 9'b10010101;
				8'b1100101: c <= 9'b101010000;
				8'b1111110: c <= 9'b11101001;
				8'b1111100: c <= 9'b100011010;
				8'b1010110: c <= 9'b111011100;
				8'b110010: c <= 9'b1001110;
				8'b1101101: c <= 9'b111110000;
				8'b100011: c <= 9'b110110011;
				8'b1110101: c <= 9'b1010110;
				8'b1111101: c <= 9'b111111001;
				8'b101001: c <= 9'b1111100;
				8'b1010010: c <= 9'b11111101;
				8'b1011000: c <= 9'b101000;
				8'b101110: c <= 9'b101111111;
				8'b1000001: c <= 9'b110101;
				default: c <= 9'b0;
			endcase
			9'b100001111 : case(di)
				8'b1000011: c <= 9'b110110011;
				8'b101000: c <= 9'b110100000;
				8'b111010: c <= 9'b101011101;
				8'b110110: c <= 9'b100101;
				8'b1100100: c <= 9'b11100111;
				8'b1000000: c <= 9'b100101111;
				8'b1110110: c <= 9'b10011100;
				8'b100101: c <= 9'b110010001;
				8'b101111: c <= 9'b101111111;
				8'b100110: c <= 9'b110111001;
				8'b1100011: c <= 9'b11111;
				8'b1001000: c <= 9'b100001001;
				8'b111000: c <= 9'b11000111;
				8'b110001: c <= 9'b100110111;
				8'b1010111: c <= 9'b111011100;
				8'b1001110: c <= 9'b1001000;
				8'b1101010: c <= 9'b111000011;
				8'b1001001: c <= 9'b11010000;
				8'b1100000: c <= 9'b10110011;
				8'b110111: c <= 9'b110000111;
				8'b1011101: c <= 9'b100110111;
				8'b1011011: c <= 9'b10101;
				8'b111001: c <= 9'b110100011;
				8'b1001010: c <= 9'b1001;
				8'b110011: c <= 9'b1101110;
				8'b1101100: c <= 9'b1011100;
				8'b1110111: c <= 9'b11001011;
				8'b101011: c <= 9'b10010011;
				8'b1101011: c <= 9'b100101111;
				8'b111100: c <= 9'b100010000;
				8'b1000111: c <= 9'b1111010;
				8'b1011111: c <= 9'b1011111;
				8'b1110100: c <= 9'b1101100;
				8'b101101: c <= 9'b101100100;
				8'b1010011: c <= 9'b111101100;
				8'b1100001: c <= 9'b100101;
				8'b110101: c <= 9'b111010010;
				8'b1000100: c <= 9'b10010101;
				8'b1010001: c <= 9'b100100101;
				8'b1010100: c <= 9'b1110000;
				8'b1100110: c <= 9'b101010100;
				8'b101010: c <= 9'b110;
				8'b1011110: c <= 9'b110100111;
				8'b1100111: c <= 9'b10011111;
				8'b1011010: c <= 9'b100011001;
				8'b1000010: c <= 9'b100000010;
				8'b111101: c <= 9'b111001111;
				8'b110000: c <= 9'b100110101;
				8'b111110: c <= 9'b101011101;
				8'b1100010: c <= 9'b11110111;
				8'b1110000: c <= 9'b101110011;
				8'b1101001: c <= 9'b11000100;
				8'b1110011: c <= 9'b10010111;
				8'b1001100: c <= 9'b101000100;
				8'b100001: c <= 9'b1100001;
				8'b1000110: c <= 9'b101100011;
				8'b1110010: c <= 9'b111001000;
				8'b1010000: c <= 9'b101100101;
				8'b1111010: c <= 9'b11110100;
				8'b1010101: c <= 9'b100110110;
				8'b111011: c <= 9'b10111000;
				8'b1001101: c <= 9'b1011001;
				8'b111111: c <= 9'b10101011;
				8'b1101110: c <= 9'b100101001;
				8'b1111011: c <= 9'b10110100;
				8'b1001011: c <= 9'b100101;
				8'b1101111: c <= 9'b101101010;
				8'b1101000: c <= 9'b101100011;
				8'b101100: c <= 9'b110101011;
				8'b100100: c <= 9'b11110;
				8'b1111000: c <= 9'b111111010;
				8'b1000101: c <= 9'b11100111;
				8'b1011001: c <= 9'b100011101;
				8'b110100: c <= 9'b101100000;
				8'b1111001: c <= 9'b10101111;
				8'b1110001: c <= 9'b10;
				8'b1001111: c <= 9'b100111011;
				8'b1100101: c <= 9'b111101010;
				8'b1111110: c <= 9'b100101111;
				8'b1111100: c <= 9'b11100101;
				8'b1010110: c <= 9'b110000111;
				8'b110010: c <= 9'b11111;
				8'b1101101: c <= 9'b11011101;
				8'b100011: c <= 9'b1000011;
				8'b1110101: c <= 9'b10110100;
				8'b1111101: c <= 9'b11010111;
				8'b101001: c <= 9'b101000110;
				8'b1010010: c <= 9'b100;
				8'b1011000: c <= 9'b1110;
				8'b101110: c <= 9'b100001001;
				8'b1000001: c <= 9'b110101011;
				default: c <= 9'b0;
			endcase
			9'b100001 : case(di)
				8'b1000011: c <= 9'b11101;
				8'b101000: c <= 9'b1111101;
				8'b111010: c <= 9'b111111110;
				8'b110110: c <= 9'b101101101;
				8'b1100100: c <= 9'b1000101;
				8'b1000000: c <= 9'b1001;
				8'b1110110: c <= 9'b11000001;
				8'b100101: c <= 9'b11101;
				8'b101111: c <= 9'b10101101;
				8'b100110: c <= 9'b1001001;
				8'b1100011: c <= 9'b100111010;
				8'b1001000: c <= 9'b110011000;
				8'b111000: c <= 9'b1000110;
				8'b110001: c <= 9'b111111001;
				8'b1010111: c <= 9'b110110;
				8'b1001110: c <= 9'b1011111;
				8'b1101010: c <= 9'b101110011;
				8'b1001001: c <= 9'b100110000;
				8'b1100000: c <= 9'b111001001;
				8'b110111: c <= 9'b101011001;
				8'b1011101: c <= 9'b1110000;
				8'b1011011: c <= 9'b110000;
				8'b111001: c <= 9'b100000010;
				8'b1001010: c <= 9'b11101111;
				8'b110011: c <= 9'b11001;
				8'b1101100: c <= 9'b101100110;
				8'b1110111: c <= 9'b101101100;
				8'b101011: c <= 9'b110000000;
				8'b1101011: c <= 9'b101010010;
				8'b111100: c <= 9'b111100000;
				8'b1000111: c <= 9'b111000;
				8'b1011111: c <= 9'b111010010;
				8'b1110100: c <= 9'b1111011;
				8'b101101: c <= 9'b100100;
				8'b1010011: c <= 9'b101001;
				8'b1100001: c <= 9'b1101110;
				8'b110101: c <= 9'b100101110;
				8'b1000100: c <= 9'b1111001;
				8'b1010001: c <= 9'b10110011;
				8'b1010100: c <= 9'b101001110;
				8'b1100110: c <= 9'b100000111;
				8'b101010: c <= 9'b1100101;
				8'b1011110: c <= 9'b100111;
				8'b1100111: c <= 9'b110110;
				8'b1011010: c <= 9'b10100;
				8'b1000010: c <= 9'b11001100;
				8'b111101: c <= 9'b110001100;
				8'b110000: c <= 9'b1001100;
				8'b111110: c <= 9'b1101110;
				8'b1100010: c <= 9'b1000101;
				8'b1110000: c <= 9'b110010001;
				8'b1101001: c <= 9'b11000001;
				8'b1110011: c <= 9'b10000010;
				8'b1001100: c <= 9'b110010011;
				8'b100001: c <= 9'b111001011;
				8'b1000110: c <= 9'b101010101;
				8'b1110010: c <= 9'b110011000;
				8'b1010000: c <= 9'b101110001;
				8'b1111010: c <= 9'b101100001;
				8'b1010101: c <= 9'b101000;
				8'b111011: c <= 9'b111010110;
				8'b1001101: c <= 9'b111111011;
				8'b111111: c <= 9'b111111101;
				8'b1101110: c <= 9'b110110000;
				8'b1111011: c <= 9'b101100111;
				8'b1001011: c <= 9'b11000;
				8'b1101111: c <= 9'b11111100;
				8'b1101000: c <= 9'b10100101;
				8'b101100: c <= 9'b111011010;
				8'b100100: c <= 9'b1011000;
				8'b1111000: c <= 9'b10111;
				8'b1000101: c <= 9'b10110111;
				8'b1011001: c <= 9'b111100101;
				8'b110100: c <= 9'b111000010;
				8'b1111001: c <= 9'b10010;
				8'b1110001: c <= 9'b100111101;
				8'b1001111: c <= 9'b11111001;
				8'b1100101: c <= 9'b10011;
				8'b1111110: c <= 9'b1110;
				8'b1111100: c <= 9'b101001100;
				8'b1010110: c <= 9'b110110;
				8'b110010: c <= 9'b11001;
				8'b1101101: c <= 9'b1101010;
				8'b100011: c <= 9'b11010001;
				8'b1110101: c <= 9'b100001101;
				8'b1111101: c <= 9'b10001110;
				8'b101001: c <= 9'b11110;
				8'b1010010: c <= 9'b1001001;
				8'b1011000: c <= 9'b100110110;
				8'b101110: c <= 9'b100011100;
				8'b1000001: c <= 9'b100001;
				default: c <= 9'b0;
			endcase
			9'b100010010 : case(di)
				8'b1000011: c <= 9'b110100000;
				8'b101000: c <= 9'b100001001;
				8'b111010: c <= 9'b110101100;
				8'b110110: c <= 9'b11000000;
				8'b1100100: c <= 9'b100111111;
				8'b1000000: c <= 9'b101001111;
				8'b1110110: c <= 9'b101111000;
				8'b100101: c <= 9'b100000010;
				8'b101111: c <= 9'b10011111;
				8'b100110: c <= 9'b110100011;
				8'b1100011: c <= 9'b111001101;
				8'b1001000: c <= 9'b111001;
				8'b111000: c <= 9'b10110101;
				8'b110001: c <= 9'b110110000;
				8'b1010111: c <= 9'b100101001;
				8'b1001110: c <= 9'b100110000;
				8'b1101010: c <= 9'b10010101;
				8'b1001001: c <= 9'b111011;
				8'b1100000: c <= 9'b110110000;
				8'b110111: c <= 9'b100100000;
				8'b1011101: c <= 9'b100011000;
				8'b1011011: c <= 9'b111110110;
				8'b111001: c <= 9'b1000010;
				8'b1001010: c <= 9'b11110101;
				8'b110011: c <= 9'b101111110;
				8'b1101100: c <= 9'b101010011;
				8'b1110111: c <= 9'b101011110;
				8'b101011: c <= 9'b10110;
				8'b1101011: c <= 9'b111000111;
				8'b111100: c <= 9'b111000100;
				8'b1000111: c <= 9'b110000;
				8'b1011111: c <= 9'b100110101;
				8'b1110100: c <= 9'b11110000;
				8'b101101: c <= 9'b11;
				8'b1010011: c <= 9'b111001001;
				8'b1100001: c <= 9'b11100011;
				8'b110101: c <= 9'b11100001;
				8'b1000100: c <= 9'b100100110;
				8'b1010001: c <= 9'b10000011;
				8'b1010100: c <= 9'b101101010;
				8'b1100110: c <= 9'b1100011;
				8'b101010: c <= 9'b101000011;
				8'b1011110: c <= 9'b100110111;
				8'b1100111: c <= 9'b111111011;
				8'b1011010: c <= 9'b111100110;
				8'b1000010: c <= 9'b1101010;
				8'b111101: c <= 9'b11110010;
				8'b110000: c <= 9'b11100010;
				8'b111110: c <= 9'b101111110;
				8'b1100010: c <= 9'b1010101;
				8'b1110000: c <= 9'b11001000;
				8'b1101001: c <= 9'b111000;
				8'b1110011: c <= 9'b11001100;
				8'b1001100: c <= 9'b11010;
				8'b100001: c <= 9'b110010;
				8'b1000110: c <= 9'b111110011;
				8'b1110010: c <= 9'b1010111;
				8'b1010000: c <= 9'b10111;
				8'b1111010: c <= 9'b100011000;
				8'b1010101: c <= 9'b111101101;
				8'b111011: c <= 9'b100111110;
				8'b1001101: c <= 9'b100101001;
				8'b111111: c <= 9'b100011011;
				8'b1101110: c <= 9'b11111001;
				8'b1111011: c <= 9'b100110111;
				8'b1001011: c <= 9'b10011;
				8'b1101111: c <= 9'b1;
				8'b1101000: c <= 9'b1011011;
				8'b101100: c <= 9'b11110111;
				8'b100100: c <= 9'b10110110;
				8'b1111000: c <= 9'b101010;
				8'b1000101: c <= 9'b101000001;
				8'b1011001: c <= 9'b110001;
				8'b110100: c <= 9'b1111000;
				8'b1111001: c <= 9'b101110111;
				8'b1110001: c <= 9'b1111110;
				8'b1001111: c <= 9'b11110111;
				8'b1100101: c <= 9'b111110000;
				8'b1111110: c <= 9'b1101001;
				8'b1111100: c <= 9'b10100010;
				8'b1010110: c <= 9'b111100110;
				8'b110010: c <= 9'b11111010;
				8'b1101101: c <= 9'b100011101;
				8'b100011: c <= 9'b100000001;
				8'b1110101: c <= 9'b101110111;
				8'b1111101: c <= 9'b10101010;
				8'b101001: c <= 9'b110101010;
				8'b1010010: c <= 9'b1100001;
				8'b1011000: c <= 9'b110000011;
				8'b101110: c <= 9'b101101100;
				8'b1000001: c <= 9'b1001100;
				default: c <= 9'b0;
			endcase
			9'b100110101 : case(di)
				8'b1000011: c <= 9'b10110001;
				8'b101000: c <= 9'b1010110;
				8'b111010: c <= 9'b10010110;
				8'b110110: c <= 9'b11100100;
				8'b1100100: c <= 9'b110011110;
				8'b1000000: c <= 9'b101101101;
				8'b1110110: c <= 9'b11100011;
				8'b100101: c <= 9'b11111110;
				8'b101111: c <= 9'b101011111;
				8'b100110: c <= 9'b1110100;
				8'b1100011: c <= 9'b111001001;
				8'b1001000: c <= 9'b110010010;
				8'b111000: c <= 9'b11000001;
				8'b110001: c <= 9'b110010110;
				8'b1010111: c <= 9'b101100110;
				8'b1001110: c <= 9'b11101111;
				8'b1101010: c <= 9'b110;
				8'b1001001: c <= 9'b11101100;
				8'b1100000: c <= 9'b11100101;
				8'b110111: c <= 9'b110001011;
				8'b1011101: c <= 9'b100001010;
				8'b1011011: c <= 9'b111111010;
				8'b111001: c <= 9'b101100111;
				8'b1001010: c <= 9'b111101001;
				8'b110011: c <= 9'b101101011;
				8'b1101100: c <= 9'b11001100;
				8'b1110111: c <= 9'b1111100;
				8'b101011: c <= 9'b11101001;
				8'b1101011: c <= 9'b100111010;
				8'b111100: c <= 9'b1100011;
				8'b1000111: c <= 9'b100101011;
				8'b1011111: c <= 9'b100010010;
				8'b1110100: c <= 9'b1001001;
				8'b101101: c <= 9'b101010101;
				8'b1010011: c <= 9'b10010101;
				8'b1100001: c <= 9'b10000001;
				8'b110101: c <= 9'b100001;
				8'b1000100: c <= 9'b111001101;
				8'b1010001: c <= 9'b11100110;
				8'b1010100: c <= 9'b110111010;
				8'b1100110: c <= 9'b100110100;
				8'b101010: c <= 9'b100101;
				8'b1011110: c <= 9'b101001110;
				8'b1100111: c <= 9'b110110100;
				8'b1011010: c <= 9'b110000;
				8'b1000010: c <= 9'b10001001;
				8'b111101: c <= 9'b11101111;
				8'b110000: c <= 9'b11100100;
				8'b111110: c <= 9'b1100000;
				8'b1100010: c <= 9'b110111;
				8'b1110000: c <= 9'b110001001;
				8'b1101001: c <= 9'b110011000;
				8'b1110011: c <= 9'b111010100;
				8'b1001100: c <= 9'b110111010;
				8'b100001: c <= 9'b1000;
				8'b1000110: c <= 9'b101010;
				8'b1110010: c <= 9'b1111011;
				8'b1010000: c <= 9'b10000011;
				8'b1111010: c <= 9'b10111000;
				8'b1010101: c <= 9'b111111011;
				8'b111011: c <= 9'b110001001;
				8'b1001101: c <= 9'b11011010;
				8'b111111: c <= 9'b10000011;
				8'b1101110: c <= 9'b111000111;
				8'b1111011: c <= 9'b11001100;
				8'b1001011: c <= 9'b10100110;
				8'b1101111: c <= 9'b10001101;
				8'b1101000: c <= 9'b10101000;
				8'b101100: c <= 9'b11010010;
				8'b100100: c <= 9'b100110010;
				8'b1111000: c <= 9'b11100011;
				8'b1000101: c <= 9'b111110011;
				8'b1011001: c <= 9'b110110101;
				8'b110100: c <= 9'b111101110;
				8'b1111001: c <= 9'b100110;
				8'b1110001: c <= 9'b110011010;
				8'b1001111: c <= 9'b1110111;
				8'b1100101: c <= 9'b10110111;
				8'b1111110: c <= 9'b100111010;
				8'b1111100: c <= 9'b1000111;
				8'b1010110: c <= 9'b100001101;
				8'b110010: c <= 9'b1010001;
				8'b1101101: c <= 9'b10100;
				8'b100011: c <= 9'b111010001;
				8'b1110101: c <= 9'b100001001;
				8'b1111101: c <= 9'b101100100;
				8'b101001: c <= 9'b101100000;
				8'b1010010: c <= 9'b111101;
				8'b1011000: c <= 9'b10111000;
				8'b101110: c <= 9'b100101000;
				8'b1000001: c <= 9'b10100000;
				default: c <= 9'b0;
			endcase
			9'b1110011 : case(di)
				8'b1000011: c <= 9'b100010;
				8'b101000: c <= 9'b101100000;
				8'b111010: c <= 9'b1101001;
				8'b110110: c <= 9'b1110010;
				8'b1100100: c <= 9'b111000111;
				8'b1000000: c <= 9'b111011001;
				8'b1110110: c <= 9'b100100010;
				8'b100101: c <= 9'b100011001;
				8'b101111: c <= 9'b101110100;
				8'b100110: c <= 9'b10110101;
				8'b1100011: c <= 9'b1001000;
				8'b1001000: c <= 9'b11110010;
				8'b111000: c <= 9'b11001100;
				8'b110001: c <= 9'b101100101;
				8'b1010111: c <= 9'b100111010;
				8'b1001110: c <= 9'b10001000;
				8'b1101010: c <= 9'b111100;
				8'b1001001: c <= 9'b101110001;
				8'b1100000: c <= 9'b111100000;
				8'b110111: c <= 9'b1100110;
				8'b1011101: c <= 9'b101110011;
				8'b1011011: c <= 9'b11000000;
				8'b111001: c <= 9'b11010010;
				8'b1001010: c <= 9'b11001110;
				8'b110011: c <= 9'b101111000;
				8'b1101100: c <= 9'b100000000;
				8'b1110111: c <= 9'b1101100;
				8'b101011: c <= 9'b100101111;
				8'b1101011: c <= 9'b10111001;
				8'b111100: c <= 9'b100100101;
				8'b1000111: c <= 9'b101010;
				8'b1011111: c <= 9'b110100100;
				8'b1110100: c <= 9'b1100100;
				8'b101101: c <= 9'b101010011;
				8'b1010011: c <= 9'b1001110;
				8'b1100001: c <= 9'b100110;
				8'b110101: c <= 9'b1100101;
				8'b1000100: c <= 9'b11110011;
				8'b1010001: c <= 9'b1100111;
				8'b1010100: c <= 9'b11011100;
				8'b1100110: c <= 9'b10001100;
				8'b101010: c <= 9'b110111000;
				8'b1011110: c <= 9'b111101101;
				8'b1100111: c <= 9'b11110101;
				8'b1011010: c <= 9'b100111;
				8'b1000010: c <= 9'b110010110;
				8'b111101: c <= 9'b110001100;
				8'b110000: c <= 9'b1110011;
				8'b111110: c <= 9'b1001111;
				8'b1100010: c <= 9'b111010001;
				8'b1110000: c <= 9'b110110101;
				8'b1101001: c <= 9'b111111101;
				8'b1110011: c <= 9'b111101;
				8'b1001100: c <= 9'b111001100;
				8'b100001: c <= 9'b10000111;
				8'b1000110: c <= 9'b111000110;
				8'b1110010: c <= 9'b110011111;
				8'b1010000: c <= 9'b11011;
				8'b1111010: c <= 9'b111;
				8'b1010101: c <= 9'b10101110;
				8'b111011: c <= 9'b111010111;
				8'b1001101: c <= 9'b110110111;
				8'b111111: c <= 9'b101011101;
				8'b1101110: c <= 9'b10001011;
				8'b1111011: c <= 9'b100110011;
				8'b1001011: c <= 9'b11011011;
				8'b1101111: c <= 9'b111011;
				8'b1101000: c <= 9'b111111010;
				8'b101100: c <= 9'b110001;
				8'b100100: c <= 9'b111100111;
				8'b1111000: c <= 9'b101010000;
				8'b1000101: c <= 9'b1100001;
				8'b1011001: c <= 9'b10011011;
				8'b110100: c <= 9'b11101000;
				8'b1111001: c <= 9'b101100;
				8'b1110001: c <= 9'b100101010;
				8'b1001111: c <= 9'b10101101;
				8'b1100101: c <= 9'b11011101;
				8'b1111110: c <= 9'b11110010;
				8'b1111100: c <= 9'b11011010;
				8'b1010110: c <= 9'b111101010;
				8'b110010: c <= 9'b1101100;
				8'b1101101: c <= 9'b101110;
				8'b100011: c <= 9'b1010000;
				8'b1110101: c <= 9'b11000100;
				8'b1111101: c <= 9'b11000001;
				8'b101001: c <= 9'b101011;
				8'b1010010: c <= 9'b100110100;
				8'b1011000: c <= 9'b11000001;
				8'b101110: c <= 9'b101011110;
				8'b1000001: c <= 9'b111110011;
				default: c <= 9'b0;
			endcase
			9'b10110100 : case(di)
				8'b1000011: c <= 9'b101101;
				8'b101000: c <= 9'b111101111;
				8'b111010: c <= 9'b11011101;
				8'b110110: c <= 9'b10101010;
				8'b1100100: c <= 9'b111000011;
				8'b1000000: c <= 9'b1110001;
				8'b1110110: c <= 9'b11001111;
				8'b100101: c <= 9'b11101001;
				8'b101111: c <= 9'b10011101;
				8'b100110: c <= 9'b111011;
				8'b1100011: c <= 9'b11011000;
				8'b1001000: c <= 9'b11111010;
				8'b111000: c <= 9'b1101001;
				8'b110001: c <= 9'b10000111;
				8'b1010111: c <= 9'b111111001;
				8'b1001110: c <= 9'b111100101;
				8'b1101010: c <= 9'b10011010;
				8'b1001001: c <= 9'b11111;
				8'b1100000: c <= 9'b110101111;
				8'b110111: c <= 9'b11001011;
				8'b1011101: c <= 9'b100010010;
				8'b1011011: c <= 9'b100001111;
				8'b111001: c <= 9'b100001110;
				8'b1001010: c <= 9'b11010010;
				8'b110011: c <= 9'b111100010;
				8'b1101100: c <= 9'b110101;
				8'b1110111: c <= 9'b1100000;
				8'b101011: c <= 9'b10000000;
				8'b1101011: c <= 9'b10101;
				8'b111100: c <= 9'b111000101;
				8'b1000111: c <= 9'b100000000;
				8'b1011111: c <= 9'b110011111;
				8'b1110100: c <= 9'b101010100;
				8'b101101: c <= 9'b110010010;
				8'b1010011: c <= 9'b101100001;
				8'b1100001: c <= 9'b110101010;
				8'b110101: c <= 9'b110101100;
				8'b1000100: c <= 9'b100010110;
				8'b1010001: c <= 9'b10111001;
				8'b1010100: c <= 9'b11000010;
				8'b1100110: c <= 9'b110110100;
				8'b101010: c <= 9'b10001001;
				8'b1011110: c <= 9'b110;
				8'b1100111: c <= 9'b101010010;
				8'b1011010: c <= 9'b10110111;
				8'b1000010: c <= 9'b101010000;
				8'b111101: c <= 9'b111101001;
				8'b110000: c <= 9'b11100001;
				8'b111110: c <= 9'b10111111;
				8'b1100010: c <= 9'b1010011;
				8'b1110000: c <= 9'b110101010;
				8'b1101001: c <= 9'b1011010;
				8'b1110011: c <= 9'b111;
				8'b1001100: c <= 9'b110011001;
				8'b100001: c <= 9'b101001011;
				8'b1000110: c <= 9'b111101111;
				8'b1110010: c <= 9'b11001011;
				8'b1010000: c <= 9'b111111111;
				8'b1111010: c <= 9'b111001111;
				8'b1010101: c <= 9'b100010100;
				8'b111011: c <= 9'b10010001;
				8'b1001101: c <= 9'b101110001;
				8'b111111: c <= 9'b1100110;
				8'b1101110: c <= 9'b10110011;
				8'b1111011: c <= 9'b100100;
				8'b1001011: c <= 9'b1011111;
				8'b1101111: c <= 9'b110101111;
				8'b1101000: c <= 9'b11111110;
				8'b101100: c <= 9'b101001010;
				8'b100100: c <= 9'b11100000;
				8'b1111000: c <= 9'b101111001;
				8'b1000101: c <= 9'b100000011;
				8'b1011001: c <= 9'b101011101;
				8'b110100: c <= 9'b10101110;
				8'b1111001: c <= 9'b100111000;
				8'b1110001: c <= 9'b110000010;
				8'b1001111: c <= 9'b10000010;
				8'b1100101: c <= 9'b110001010;
				8'b1111110: c <= 9'b11110110;
				8'b1111100: c <= 9'b111111010;
				8'b1010110: c <= 9'b101101101;
				8'b110010: c <= 9'b11111100;
				8'b1101101: c <= 9'b10101101;
				8'b100011: c <= 9'b100010010;
				8'b1110101: c <= 9'b111001010;
				8'b1111101: c <= 9'b100001;
				8'b101001: c <= 9'b101011010;
				8'b1010010: c <= 9'b100001001;
				8'b1011000: c <= 9'b110001101;
				8'b101110: c <= 9'b10101001;
				8'b1000001: c <= 9'b111000100;
				default: c <= 9'b0;
			endcase
			9'b11011100 : case(di)
				8'b1000011: c <= 9'b110001101;
				8'b101000: c <= 9'b100011001;
				8'b111010: c <= 9'b11000;
				8'b110110: c <= 9'b111000011;
				8'b1100100: c <= 9'b110000011;
				8'b1000000: c <= 9'b11000000;
				8'b1110110: c <= 9'b1100110;
				8'b100101: c <= 9'b100101010;
				8'b101111: c <= 9'b110100100;
				8'b100110: c <= 9'b10010100;
				8'b1100011: c <= 9'b110;
				8'b1001000: c <= 9'b111001111;
				8'b111000: c <= 9'b10010111;
				8'b110001: c <= 9'b101011111;
				8'b1010111: c <= 9'b10111111;
				8'b1001110: c <= 9'b1111111;
				8'b1101010: c <= 9'b11110010;
				8'b1001001: c <= 9'b11100;
				8'b1100000: c <= 9'b1100110;
				8'b110111: c <= 9'b110010011;
				8'b1011101: c <= 9'b100111100;
				8'b1011011: c <= 9'b100111101;
				8'b111001: c <= 9'b111001000;
				8'b1001010: c <= 9'b101101010;
				8'b110011: c <= 9'b101100110;
				8'b1101100: c <= 9'b11001011;
				8'b1110111: c <= 9'b110010101;
				8'b101011: c <= 9'b100010111;
				8'b1101011: c <= 9'b100111101;
				8'b111100: c <= 9'b10110011;
				8'b1000111: c <= 9'b100010110;
				8'b1011111: c <= 9'b100110;
				8'b1110100: c <= 9'b1011;
				8'b101101: c <= 9'b111001010;
				8'b1010011: c <= 9'b11110010;
				8'b1100001: c <= 9'b111101110;
				8'b110101: c <= 9'b10011011;
				8'b1000100: c <= 9'b100110100;
				8'b1010001: c <= 9'b100011010;
				8'b1010100: c <= 9'b1011110;
				8'b1100110: c <= 9'b110001111;
				8'b101010: c <= 9'b101110;
				8'b1011110: c <= 9'b111110011;
				8'b1100111: c <= 9'b10000111;
				8'b1011010: c <= 9'b111001000;
				8'b1000010: c <= 9'b101011000;
				8'b111101: c <= 9'b100100011;
				8'b110000: c <= 9'b10101010;
				8'b111110: c <= 9'b100101001;
				8'b1100010: c <= 9'b100111101;
				8'b1110000: c <= 9'b111101100;
				8'b1101001: c <= 9'b10011101;
				8'b1110011: c <= 9'b110100101;
				8'b1001100: c <= 9'b10110111;
				8'b100001: c <= 9'b101010010;
				8'b1000110: c <= 9'b101101000;
				8'b1110010: c <= 9'b111100001;
				8'b1010000: c <= 9'b110110100;
				8'b1111010: c <= 9'b111101100;
				8'b1010101: c <= 9'b10001011;
				8'b111011: c <= 9'b10101000;
				8'b1001101: c <= 9'b10111000;
				8'b111111: c <= 9'b11001100;
				8'b1101110: c <= 9'b101100011;
				8'b1111011: c <= 9'b10001001;
				8'b1001011: c <= 9'b11100110;
				8'b1101111: c <= 9'b11011011;
				8'b1101000: c <= 9'b111101001;
				8'b101100: c <= 9'b11111001;
				8'b100100: c <= 9'b10100111;
				8'b1111000: c <= 9'b11011110;
				8'b1000101: c <= 9'b1011100;
				8'b1011001: c <= 9'b100101100;
				8'b110100: c <= 9'b1000110;
				8'b1111001: c <= 9'b101110011;
				8'b1110001: c <= 9'b101001010;
				8'b1001111: c <= 9'b11111101;
				8'b1100101: c <= 9'b1101000;
				8'b1111110: c <= 9'b1101111;
				8'b1111100: c <= 9'b100011101;
				8'b1010110: c <= 9'b100110110;
				8'b110010: c <= 9'b101010;
				8'b1101101: c <= 9'b100010000;
				8'b100011: c <= 9'b101111010;
				8'b1110101: c <= 9'b11101000;
				8'b1111101: c <= 9'b11111101;
				8'b101001: c <= 9'b110101111;
				8'b1010010: c <= 9'b100000100;
				8'b1011000: c <= 9'b1111;
				8'b101110: c <= 9'b10110110;
				8'b1000001: c <= 9'b100000011;
				default: c <= 9'b0;
			endcase
			9'b111011110 : case(di)
				8'b1000011: c <= 9'b10100011;
				8'b101000: c <= 9'b110110101;
				8'b111010: c <= 9'b101101010;
				8'b110110: c <= 9'b111001000;
				8'b1100100: c <= 9'b100010010;
				8'b1000000: c <= 9'b110101001;
				8'b1110110: c <= 9'b110100000;
				8'b100101: c <= 9'b101010001;
				8'b101111: c <= 9'b101111001;
				8'b100110: c <= 9'b110101011;
				8'b1100011: c <= 9'b1010110;
				8'b1001000: c <= 9'b110110100;
				8'b111000: c <= 9'b100001011;
				8'b110001: c <= 9'b100101010;
				8'b1010111: c <= 9'b111100101;
				8'b1001110: c <= 9'b110111110;
				8'b1101010: c <= 9'b111000101;
				8'b1001001: c <= 9'b111110110;
				8'b1100000: c <= 9'b100110101;
				8'b110111: c <= 9'b111111011;
				8'b1011101: c <= 9'b1110000;
				8'b1011011: c <= 9'b11110011;
				8'b111001: c <= 9'b11101100;
				8'b1001010: c <= 9'b110000110;
				8'b110011: c <= 9'b1001111;
				8'b1101100: c <= 9'b11000110;
				8'b1110111: c <= 9'b110011010;
				8'b101011: c <= 9'b101000001;
				8'b1101011: c <= 9'b1011111;
				8'b111100: c <= 9'b11011011;
				8'b1000111: c <= 9'b101000111;
				8'b1011111: c <= 9'b110101110;
				8'b1110100: c <= 9'b100011001;
				8'b101101: c <= 9'b100111010;
				8'b1010011: c <= 9'b111111111;
				8'b1100001: c <= 9'b10000111;
				8'b110101: c <= 9'b100011011;
				8'b1000100: c <= 9'b11101100;
				8'b1010001: c <= 9'b101010111;
				8'b1010100: c <= 9'b100010010;
				8'b1100110: c <= 9'b110001001;
				8'b101010: c <= 9'b110010100;
				8'b1011110: c <= 9'b1111111;
				8'b1100111: c <= 9'b110000010;
				8'b1011010: c <= 9'b101110;
				8'b1000010: c <= 9'b1100101;
				8'b111101: c <= 9'b11100111;
				8'b110000: c <= 9'b11100101;
				8'b111110: c <= 9'b110101101;
				8'b1100010: c <= 9'b111101110;
				8'b1110000: c <= 9'b11110111;
				8'b1101001: c <= 9'b111010010;
				8'b1110011: c <= 9'b101100100;
				8'b1001100: c <= 9'b111010000;
				8'b100001: c <= 9'b111011111;
				8'b1000110: c <= 9'b1100100;
				8'b1110010: c <= 9'b1101000;
				8'b1010000: c <= 9'b10;
				8'b1111010: c <= 9'b110001100;
				8'b1010101: c <= 9'b10011000;
				8'b111011: c <= 9'b110010011;
				8'b1001101: c <= 9'b100110011;
				8'b111111: c <= 9'b110010101;
				8'b1101110: c <= 9'b1101001;
				8'b1111011: c <= 9'b101101;
				8'b1001011: c <= 9'b100011101;
				8'b1101111: c <= 9'b111110001;
				8'b1101000: c <= 9'b101101011;
				8'b101100: c <= 9'b1110011;
				8'b100100: c <= 9'b110100010;
				8'b1111000: c <= 9'b110100110;
				8'b1000101: c <= 9'b100010100;
				8'b1011001: c <= 9'b111101100;
				8'b110100: c <= 9'b100111011;
				8'b1111001: c <= 9'b1011110;
				8'b1110001: c <= 9'b111110101;
				8'b1001111: c <= 9'b101010101;
				8'b1100101: c <= 9'b11101111;
				8'b1111110: c <= 9'b100110101;
				8'b1111100: c <= 9'b10011100;
				8'b1010110: c <= 9'b110111011;
				8'b110010: c <= 9'b110000;
				8'b1101101: c <= 9'b1000101;
				8'b100011: c <= 9'b111100000;
				8'b1110101: c <= 9'b1100;
				8'b1111101: c <= 9'b1000111;
				8'b101001: c <= 9'b11100010;
				8'b1010010: c <= 9'b1101100;
				8'b1011000: c <= 9'b100100;
				8'b101110: c <= 9'b11010011;
				8'b1000001: c <= 9'b111111011;
				default: c <= 9'b0;
			endcase
			9'b1110001 : case(di)
				8'b1000011: c <= 9'b10101100;
				8'b101000: c <= 9'b1100101;
				8'b111010: c <= 9'b11001000;
				8'b110110: c <= 9'b1001111;
				8'b1100100: c <= 9'b10010111;
				8'b1000000: c <= 9'b111100001;
				8'b1110110: c <= 9'b101011001;
				8'b100101: c <= 9'b110001;
				8'b101111: c <= 9'b111000110;
				8'b100110: c <= 9'b1010110;
				8'b1100011: c <= 9'b110111100;
				8'b1001000: c <= 9'b10100110;
				8'b111000: c <= 9'b111011011;
				8'b110001: c <= 9'b1110000;
				8'b1010111: c <= 9'b110101101;
				8'b1001110: c <= 9'b101101110;
				8'b1101010: c <= 9'b101101001;
				8'b1001001: c <= 9'b110000101;
				8'b1100000: c <= 9'b10000111;
				8'b110111: c <= 9'b1101111;
				8'b1011101: c <= 9'b101101011;
				8'b1011011: c <= 9'b110110000;
				8'b111001: c <= 9'b110000110;
				8'b1001010: c <= 9'b111010100;
				8'b110011: c <= 9'b100101001;
				8'b1101100: c <= 9'b10010001;
				8'b1110111: c <= 9'b11010101;
				8'b101011: c <= 9'b100100010;
				8'b1101011: c <= 9'b1101110;
				8'b111100: c <= 9'b110100010;
				8'b1000111: c <= 9'b10111111;
				8'b1011111: c <= 9'b110000;
				8'b1110100: c <= 9'b1100110;
				8'b101101: c <= 9'b100101010;
				8'b1010011: c <= 9'b11110000;
				8'b1100001: c <= 9'b101001011;
				8'b110101: c <= 9'b101000010;
				8'b1000100: c <= 9'b111011100;
				8'b1010001: c <= 9'b11110001;
				8'b1010100: c <= 9'b111011111;
				8'b1100110: c <= 9'b100100010;
				8'b101010: c <= 9'b110100100;
				8'b1011110: c <= 9'b10101110;
				8'b1100111: c <= 9'b100010000;
				8'b1011010: c <= 9'b100100011;
				8'b1000010: c <= 9'b1001111;
				8'b111101: c <= 9'b110000001;
				8'b110000: c <= 9'b11110;
				8'b111110: c <= 9'b100110101;
				8'b1100010: c <= 9'b110000110;
				8'b1110000: c <= 9'b101111111;
				8'b1101001: c <= 9'b111000;
				8'b1110011: c <= 9'b11;
				8'b1001100: c <= 9'b11101011;
				8'b100001: c <= 9'b110010;
				8'b1000110: c <= 9'b111100;
				8'b1110010: c <= 9'b1100011;
				8'b1010000: c <= 9'b101111010;
				8'b1111010: c <= 9'b1100011;
				8'b1010101: c <= 9'b110000111;
				8'b111011: c <= 9'b11000010;
				8'b1001101: c <= 9'b110010110;
				8'b111111: c <= 9'b10111110;
				8'b1101110: c <= 9'b101011001;
				8'b1111011: c <= 9'b1011010;
				8'b1001011: c <= 9'b110;
				8'b1101111: c <= 9'b110111110;
				8'b1101000: c <= 9'b101011010;
				8'b101100: c <= 9'b11001;
				8'b100100: c <= 9'b10110;
				8'b1111000: c <= 9'b111011001;
				8'b1000101: c <= 9'b1010010;
				8'b1011001: c <= 9'b111100111;
				8'b110100: c <= 9'b100010001;
				8'b1111001: c <= 9'b110001111;
				8'b1110001: c <= 9'b1101111;
				8'b1001111: c <= 9'b10101110;
				8'b1100101: c <= 9'b11101100;
				8'b1111110: c <= 9'b100101000;
				8'b1111100: c <= 9'b111000110;
				8'b1010110: c <= 9'b110001011;
				8'b110010: c <= 9'b11001111;
				8'b1101101: c <= 9'b10110100;
				8'b100011: c <= 9'b100101;
				8'b1110101: c <= 9'b110011001;
				8'b1111101: c <= 9'b100110011;
				8'b101001: c <= 9'b110101;
				8'b1010010: c <= 9'b1000101;
				8'b1011000: c <= 9'b100001100;
				8'b101110: c <= 9'b10011001;
				8'b1000001: c <= 9'b101101110;
				default: c <= 9'b0;
			endcase
			9'b101000 : case(di)
				8'b1000011: c <= 9'b1110001;
				8'b101000: c <= 9'b111110101;
				8'b111010: c <= 9'b110111001;
				8'b110110: c <= 9'b11011001;
				8'b1100100: c <= 9'b101111010;
				8'b1000000: c <= 9'b100011100;
				8'b1110110: c <= 9'b11110011;
				8'b100101: c <= 9'b100100010;
				8'b101111: c <= 9'b110011100;
				8'b100110: c <= 9'b100100110;
				8'b1100011: c <= 9'b10100100;
				8'b1001000: c <= 9'b1001000;
				8'b111000: c <= 9'b11110000;
				8'b110001: c <= 9'b11000100;
				8'b1010111: c <= 9'b111010100;
				8'b1001110: c <= 9'b1010011;
				8'b1101010: c <= 9'b1100;
				8'b1001001: c <= 9'b100001010;
				8'b1100000: c <= 9'b101010011;
				8'b110111: c <= 9'b110011010;
				8'b1011101: c <= 9'b11111010;
				8'b1011011: c <= 9'b110100100;
				8'b111001: c <= 9'b101101100;
				8'b1001010: c <= 9'b110101001;
				8'b110011: c <= 9'b10110;
				8'b1101100: c <= 9'b101000;
				8'b1110111: c <= 9'b100010011;
				8'b101011: c <= 9'b101000011;
				8'b1101011: c <= 9'b101110000;
				8'b111100: c <= 9'b10001000;
				8'b1000111: c <= 9'b100010010;
				8'b1011111: c <= 9'b10010100;
				8'b1110100: c <= 9'b110101111;
				8'b101101: c <= 9'b100000101;
				8'b1010011: c <= 9'b11000;
				8'b1100001: c <= 9'b11110010;
				8'b110101: c <= 9'b11001110;
				8'b1000100: c <= 9'b10101101;
				8'b1010001: c <= 9'b10111000;
				8'b1010100: c <= 9'b1100111;
				8'b1100110: c <= 9'b110001111;
				8'b101010: c <= 9'b11001010;
				8'b1011110: c <= 9'b110000001;
				8'b1100111: c <= 9'b110100100;
				8'b1011010: c <= 9'b1111110;
				8'b1000010: c <= 9'b111001000;
				8'b111101: c <= 9'b110111111;
				8'b110000: c <= 9'b10111;
				8'b111110: c <= 9'b100110111;
				8'b1100010: c <= 9'b1111100;
				8'b1110000: c <= 9'b101011001;
				8'b1101001: c <= 9'b100011011;
				8'b1110011: c <= 9'b10011101;
				8'b1001100: c <= 9'b111111101;
				8'b100001: c <= 9'b1001110;
				8'b1000110: c <= 9'b10000001;
				8'b1110010: c <= 9'b100000101;
				8'b1010000: c <= 9'b11000100;
				8'b1111010: c <= 9'b10011010;
				8'b1010101: c <= 9'b1;
				8'b111011: c <= 9'b1111110;
				8'b1001101: c <= 9'b100101111;
				8'b111111: c <= 9'b10000011;
				8'b1101110: c <= 9'b11111110;
				8'b1111011: c <= 9'b110010111;
				8'b1001011: c <= 9'b101111000;
				8'b1101111: c <= 9'b110011011;
				8'b1101000: c <= 9'b1100100;
				8'b101100: c <= 9'b11010001;
				8'b100100: c <= 9'b110000101;
				8'b1111000: c <= 9'b1101001;
				8'b1000101: c <= 9'b110100110;
				8'b1011001: c <= 9'b10011001;
				8'b110100: c <= 9'b110110;
				8'b1111001: c <= 9'b11111010;
				8'b1110001: c <= 9'b101011010;
				8'b1001111: c <= 9'b100100101;
				8'b1100101: c <= 9'b10001011;
				8'b1111110: c <= 9'b10101101;
				8'b1111100: c <= 9'b111111111;
				8'b1010110: c <= 9'b101011001;
				8'b110010: c <= 9'b110100000;
				8'b1101101: c <= 9'b1001011;
				8'b100011: c <= 9'b10011001;
				8'b1110101: c <= 9'b110001110;
				8'b1111101: c <= 9'b110000011;
				8'b101001: c <= 9'b11100;
				8'b1010010: c <= 9'b110011001;
				8'b1011000: c <= 9'b10101;
				8'b101110: c <= 9'b11110011;
				8'b1000001: c <= 9'b1111100;
				default: c <= 9'b0;
			endcase
			9'b10010110 : case(di)
				8'b1000011: c <= 9'b101000011;
				8'b101000: c <= 9'b100111100;
				8'b111010: c <= 9'b110001000;
				8'b110110: c <= 9'b110000011;
				8'b1100100: c <= 9'b11111110;
				8'b1000000: c <= 9'b101111000;
				8'b1110110: c <= 9'b10001100;
				8'b100101: c <= 9'b11100111;
				8'b101111: c <= 9'b101010001;
				8'b100110: c <= 9'b111011110;
				8'b1100011: c <= 9'b10101011;
				8'b1001000: c <= 9'b110111001;
				8'b111000: c <= 9'b110010;
				8'b110001: c <= 9'b100000011;
				8'b1010111: c <= 9'b1011001;
				8'b1001110: c <= 9'b11000010;
				8'b1101010: c <= 9'b1110111;
				8'b1001001: c <= 9'b101110001;
				8'b1100000: c <= 9'b1100110;
				8'b110111: c <= 9'b110010111;
				8'b1011101: c <= 9'b111010000;
				8'b1011011: c <= 9'b1110001;
				8'b111001: c <= 9'b11001101;
				8'b1001010: c <= 9'b1010000;
				8'b110011: c <= 9'b11101100;
				8'b1101100: c <= 9'b10101111;
				8'b1110111: c <= 9'b1100100;
				8'b101011: c <= 9'b100001101;
				8'b1101011: c <= 9'b101011;
				8'b111100: c <= 9'b11100001;
				8'b1000111: c <= 9'b11100000;
				8'b1011111: c <= 9'b10001111;
				8'b1110100: c <= 9'b101001;
				8'b101101: c <= 9'b100010000;
				8'b1010011: c <= 9'b1001;
				8'b1100001: c <= 9'b111101001;
				8'b110101: c <= 9'b11111101;
				8'b1000100: c <= 9'b101001111;
				8'b1010001: c <= 9'b11000000;
				8'b1010100: c <= 9'b110110100;
				8'b1100110: c <= 9'b111010100;
				8'b101010: c <= 9'b10010100;
				8'b1011110: c <= 9'b111101101;
				8'b1100111: c <= 9'b110111001;
				8'b1011010: c <= 9'b10111011;
				8'b1000010: c <= 9'b10001001;
				8'b111101: c <= 9'b1010101;
				8'b110000: c <= 9'b11001010;
				8'b111110: c <= 9'b100100110;
				8'b1100010: c <= 9'b111110110;
				8'b1110000: c <= 9'b1011001;
				8'b1101001: c <= 9'b10010011;
				8'b1110011: c <= 9'b10101000;
				8'b1001100: c <= 9'b1011011;
				8'b100001: c <= 9'b100110010;
				8'b1000110: c <= 9'b101011111;
				8'b1110010: c <= 9'b110010001;
				8'b1010000: c <= 9'b111100111;
				8'b1111010: c <= 9'b10101;
				8'b1010101: c <= 9'b100;
				8'b111011: c <= 9'b110010010;
				8'b1001101: c <= 9'b101010011;
				8'b111111: c <= 9'b11011;
				8'b1101110: c <= 9'b111010111;
				8'b1111011: c <= 9'b100001101;
				8'b1001011: c <= 9'b10011010;
				8'b1101111: c <= 9'b10100100;
				8'b1101000: c <= 9'b110100010;
				8'b101100: c <= 9'b100001101;
				8'b100100: c <= 9'b111010111;
				8'b1111000: c <= 9'b1101;
				8'b1000101: c <= 9'b111000;
				8'b1011001: c <= 9'b100001110;
				8'b110100: c <= 9'b10011010;
				8'b1111001: c <= 9'b11101111;
				8'b1110001: c <= 9'b100010101;
				8'b1001111: c <= 9'b10100100;
				8'b1100101: c <= 9'b11000010;
				8'b1111110: c <= 9'b111010;
				8'b1111100: c <= 9'b11011101;
				8'b1010110: c <= 9'b100010100;
				8'b110010: c <= 9'b111010010;
				8'b1101101: c <= 9'b10110010;
				8'b100011: c <= 9'b111011100;
				8'b1110101: c <= 9'b101111001;
				8'b1111101: c <= 9'b101;
				8'b101001: c <= 9'b101000110;
				8'b1010010: c <= 9'b1100;
				8'b1011000: c <= 9'b1111101;
				8'b101110: c <= 9'b1001011;
				8'b1000001: c <= 9'b110011010;
				default: c <= 9'b0;
			endcase
			9'b111100010 : case(di)
				8'b1000011: c <= 9'b101010000;
				8'b101000: c <= 9'b11111011;
				8'b111010: c <= 9'b10111010;
				8'b110110: c <= 9'b110001001;
				8'b1100100: c <= 9'b11000010;
				8'b1000000: c <= 9'b110110;
				8'b1110110: c <= 9'b11011011;
				8'b100101: c <= 9'b111111011;
				8'b101111: c <= 9'b10011011;
				8'b100110: c <= 9'b111011110;
				8'b1100011: c <= 9'b11010000;
				8'b1001000: c <= 9'b100110;
				8'b111000: c <= 9'b100111000;
				8'b110001: c <= 9'b111110000;
				8'b1010111: c <= 9'b101001011;
				8'b1001110: c <= 9'b10000011;
				8'b1101010: c <= 9'b111100001;
				8'b1001001: c <= 9'b110011010;
				8'b1100000: c <= 9'b111110001;
				8'b110111: c <= 9'b110010111;
				8'b1011101: c <= 9'b1101010;
				8'b1011011: c <= 9'b1011011;
				8'b111001: c <= 9'b110100;
				8'b1001010: c <= 9'b101101011;
				8'b110011: c <= 9'b110101110;
				8'b1101100: c <= 9'b111001111;
				8'b1110111: c <= 9'b101001111;
				8'b101011: c <= 9'b110110011;
				8'b1101011: c <= 9'b100110101;
				8'b111100: c <= 9'b11000100;
				8'b1000111: c <= 9'b101110111;
				8'b1011111: c <= 9'b10100100;
				8'b1110100: c <= 9'b11110100;
				8'b101101: c <= 9'b10100111;
				8'b1010011: c <= 9'b111011011;
				8'b1100001: c <= 9'b1110100;
				8'b110101: c <= 9'b100010001;
				8'b1000100: c <= 9'b1110001;
				8'b1010001: c <= 9'b101000010;
				8'b1010100: c <= 9'b100100010;
				8'b1100110: c <= 9'b11011011;
				8'b101010: c <= 9'b101101011;
				8'b1011110: c <= 9'b100111101;
				8'b1100111: c <= 9'b100011111;
				8'b1011010: c <= 9'b1000001;
				8'b1000010: c <= 9'b111100110;
				8'b111101: c <= 9'b10111101;
				8'b110000: c <= 9'b111010001;
				8'b111110: c <= 9'b110000010;
				8'b1100010: c <= 9'b100101100;
				8'b1110000: c <= 9'b110110100;
				8'b1101001: c <= 9'b100101011;
				8'b1110011: c <= 9'b11101001;
				8'b1001100: c <= 9'b110100100;
				8'b100001: c <= 9'b11000;
				8'b1000110: c <= 9'b110110100;
				8'b1110010: c <= 9'b101000;
				8'b1010000: c <= 9'b100010011;
				8'b1111010: c <= 9'b10100111;
				8'b1010101: c <= 9'b110110101;
				8'b111011: c <= 9'b1111100;
				8'b1001101: c <= 9'b111001000;
				8'b111111: c <= 9'b10101101;
				8'b1101110: c <= 9'b11010011;
				8'b1111011: c <= 9'b11000110;
				8'b1001011: c <= 9'b10001111;
				8'b1101111: c <= 9'b110000000;
				8'b1101000: c <= 9'b111101000;
				8'b101100: c <= 9'b10100;
				8'b100100: c <= 9'b1010110;
				8'b1111000: c <= 9'b100010010;
				8'b1000101: c <= 9'b100111111;
				8'b1011001: c <= 9'b10101111;
				8'b110100: c <= 9'b100110011;
				8'b1111001: c <= 9'b101010111;
				8'b1110001: c <= 9'b1010001;
				8'b1001111: c <= 9'b111000;
				8'b1100101: c <= 9'b10011101;
				8'b1111110: c <= 9'b10000000;
				8'b1111100: c <= 9'b1011000;
				8'b1010110: c <= 9'b101001010;
				8'b110010: c <= 9'b11100100;
				8'b1101101: c <= 9'b101100111;
				8'b100011: c <= 9'b110011110;
				8'b1110101: c <= 9'b100001110;
				8'b1111101: c <= 9'b101010111;
				8'b101001: c <= 9'b101010010;
				8'b1010010: c <= 9'b111111011;
				8'b1011000: c <= 9'b111100;
				8'b101110: c <= 9'b110010100;
				8'b1000001: c <= 9'b111010;
				default: c <= 9'b0;
			endcase
			9'b10101000 : case(di)
				8'b1000011: c <= 9'b110011011;
				8'b101000: c <= 9'b1000110;
				8'b111010: c <= 9'b111100111;
				8'b110110: c <= 9'b100101011;
				8'b1100100: c <= 9'b10110110;
				8'b1000000: c <= 9'b1100010;
				8'b1110110: c <= 9'b1110011;
				8'b100101: c <= 9'b100011011;
				8'b101111: c <= 9'b11110001;
				8'b100110: c <= 9'b11110100;
				8'b1100011: c <= 9'b110000101;
				8'b1001000: c <= 9'b110001;
				8'b111000: c <= 9'b10010111;
				8'b110001: c <= 9'b101000100;
				8'b1010111: c <= 9'b111111101;
				8'b1001110: c <= 9'b11101011;
				8'b1101010: c <= 9'b111111110;
				8'b1001001: c <= 9'b11011;
				8'b1100000: c <= 9'b101;
				8'b110111: c <= 9'b10010;
				8'b1011101: c <= 9'b101101001;
				8'b1011011: c <= 9'b101010;
				8'b111001: c <= 9'b10010110;
				8'b1001010: c <= 9'b110111010;
				8'b110011: c <= 9'b101111111;
				8'b1101100: c <= 9'b11100010;
				8'b1110111: c <= 9'b10000110;
				8'b101011: c <= 9'b1100111;
				8'b1101011: c <= 9'b101100100;
				8'b111100: c <= 9'b101110101;
				8'b1000111: c <= 9'b11111011;
				8'b1011111: c <= 9'b100011111;
				8'b1110100: c <= 9'b110111111;
				8'b101101: c <= 9'b110101011;
				8'b1010011: c <= 9'b100100000;
				8'b1100001: c <= 9'b11110;
				8'b110101: c <= 9'b110010001;
				8'b1000100: c <= 9'b11101101;
				8'b1010001: c <= 9'b11011;
				8'b1010100: c <= 9'b101101010;
				8'b1100110: c <= 9'b101011;
				8'b101010: c <= 9'b11000110;
				8'b1011110: c <= 9'b111000011;
				8'b1100111: c <= 9'b110001111;
				8'b1011010: c <= 9'b100111;
				8'b1000010: c <= 9'b10001111;
				8'b111101: c <= 9'b111110011;
				8'b110000: c <= 9'b1101;
				8'b111110: c <= 9'b111100;
				8'b1100010: c <= 9'b10101110;
				8'b1110000: c <= 9'b111000110;
				8'b1101001: c <= 9'b1101000;
				8'b1110011: c <= 9'b11110101;
				8'b1001100: c <= 9'b100001111;
				8'b100001: c <= 9'b1001101;
				8'b1000110: c <= 9'b111110001;
				8'b1110010: c <= 9'b1010101;
				8'b1010000: c <= 9'b1010011;
				8'b1111010: c <= 9'b101100;
				8'b1010101: c <= 9'b1010011;
				8'b111011: c <= 9'b101010100;
				8'b1001101: c <= 9'b110011010;
				8'b111111: c <= 9'b110101100;
				8'b1101110: c <= 9'b101011000;
				8'b1111011: c <= 9'b100110110;
				8'b1001011: c <= 9'b11010001;
				8'b1101111: c <= 9'b111000;
				8'b1101000: c <= 9'b110000111;
				8'b101100: c <= 9'b101010100;
				8'b100100: c <= 9'b101101101;
				8'b1111000: c <= 9'b1101110;
				8'b1000101: c <= 9'b110011001;
				8'b1011001: c <= 9'b100111110;
				8'b110100: c <= 9'b111110011;
				8'b1111001: c <= 9'b110101;
				8'b1110001: c <= 9'b101100011;
				8'b1001111: c <= 9'b100001101;
				8'b1100101: c <= 9'b1111010;
				8'b1111110: c <= 9'b101101001;
				8'b1111100: c <= 9'b11111101;
				8'b1010110: c <= 9'b10110110;
				8'b110010: c <= 9'b110110110;
				8'b1101101: c <= 9'b1101110;
				8'b100011: c <= 9'b11011;
				8'b1110101: c <= 9'b110001011;
				8'b1111101: c <= 9'b1000001;
				8'b101001: c <= 9'b101101011;
				8'b1010010: c <= 9'b1001110;
				8'b1011000: c <= 9'b11110101;
				8'b101110: c <= 9'b100;
				8'b1000001: c <= 9'b10;
				default: c <= 9'b0;
			endcase
			9'b101010001 : case(di)
				8'b1000011: c <= 9'b10111000;
				8'b101000: c <= 9'b10101001;
				8'b111010: c <= 9'b1100100;
				8'b110110: c <= 9'b10100011;
				8'b1100100: c <= 9'b111110001;
				8'b1000000: c <= 9'b110111100;
				8'b1110110: c <= 9'b10111101;
				8'b100101: c <= 9'b1100100;
				8'b101111: c <= 9'b111010;
				8'b100110: c <= 9'b100011101;
				8'b1100011: c <= 9'b101000011;
				8'b1001000: c <= 9'b101000001;
				8'b111000: c <= 9'b10011101;
				8'b110001: c <= 9'b1000111;
				8'b1010111: c <= 9'b10111011;
				8'b1001110: c <= 9'b101011001;
				8'b1101010: c <= 9'b101001100;
				8'b1001001: c <= 9'b1101010;
				8'b1100000: c <= 9'b100000011;
				8'b110111: c <= 9'b1001100;
				8'b1011101: c <= 9'b111101101;
				8'b1011011: c <= 9'b101001011;
				8'b111001: c <= 9'b11010101;
				8'b1001010: c <= 9'b10000110;
				8'b110011: c <= 9'b100110000;
				8'b1101100: c <= 9'b1101100;
				8'b1110111: c <= 9'b110110011;
				8'b101011: c <= 9'b111110110;
				8'b1101011: c <= 9'b1011010;
				8'b111100: c <= 9'b10111010;
				8'b1000111: c <= 9'b11000100;
				8'b1011111: c <= 9'b110010110;
				8'b1110100: c <= 9'b11111110;
				8'b101101: c <= 9'b10110;
				8'b1010011: c <= 9'b110000111;
				8'b1100001: c <= 9'b111111110;
				8'b110101: c <= 9'b100110101;
				8'b1000100: c <= 9'b110001001;
				8'b1010001: c <= 9'b1111011;
				8'b1010100: c <= 9'b10110100;
				8'b1100110: c <= 9'b111001011;
				8'b101010: c <= 9'b11110011;
				8'b1011110: c <= 9'b1111000;
				8'b1100111: c <= 9'b101110011;
				8'b1011010: c <= 9'b101000011;
				8'b1000010: c <= 9'b111000011;
				8'b111101: c <= 9'b100110111;
				8'b110000: c <= 9'b11100001;
				8'b111110: c <= 9'b100100001;
				8'b1100010: c <= 9'b1010110;
				8'b1110000: c <= 9'b110110;
				8'b1101001: c <= 9'b110001100;
				8'b1110011: c <= 9'b111000111;
				8'b1001100: c <= 9'b1001;
				8'b100001: c <= 9'b111100010;
				8'b1000110: c <= 9'b101100111;
				8'b1110010: c <= 9'b101110110;
				8'b1010000: c <= 9'b101100011;
				8'b1111010: c <= 9'b11100000;
				8'b1010101: c <= 9'b100111011;
				8'b111011: c <= 9'b101010101;
				8'b1001101: c <= 9'b110000000;
				8'b111111: c <= 9'b111001111;
				8'b1101110: c <= 9'b11111;
				8'b1111011: c <= 9'b1000101;
				8'b1001011: c <= 9'b11110011;
				8'b1101111: c <= 9'b1101001;
				8'b1101000: c <= 9'b1001001;
				8'b101100: c <= 9'b111111101;
				8'b100100: c <= 9'b101110;
				8'b1111000: c <= 9'b100011011;
				8'b1000101: c <= 9'b1111100;
				8'b1011001: c <= 9'b110000001;
				8'b110100: c <= 9'b10100010;
				8'b1111001: c <= 9'b111010010;
				8'b1110001: c <= 9'b1001111;
				8'b1001111: c <= 9'b110110110;
				8'b1100101: c <= 9'b111011010;
				8'b1111110: c <= 9'b11100010;
				8'b1111100: c <= 9'b111111001;
				8'b1010110: c <= 9'b110101110;
				8'b110010: c <= 9'b1010000;
				8'b1101101: c <= 9'b110110011;
				8'b100011: c <= 9'b11001110;
				8'b1110101: c <= 9'b11001;
				8'b1111101: c <= 9'b11000100;
				8'b101001: c <= 9'b110111001;
				8'b1010010: c <= 9'b11011110;
				8'b1011000: c <= 9'b110100111;
				8'b101110: c <= 9'b11000;
				8'b1000001: c <= 9'b101110111;
				default: c <= 9'b0;
			endcase
			9'b1001111 : case(di)
				8'b1000011: c <= 9'b11010111;
				8'b101000: c <= 9'b111011110;
				8'b111010: c <= 9'b111101;
				8'b110110: c <= 9'b1100;
				8'b1100100: c <= 9'b100100010;
				8'b1000000: c <= 9'b10;
				8'b1110110: c <= 9'b100001001;
				8'b100101: c <= 9'b11000010;
				8'b101111: c <= 9'b10011011;
				8'b100110: c <= 9'b111111;
				8'b1100011: c <= 9'b110011111;
				8'b1001000: c <= 9'b101011110;
				8'b111000: c <= 9'b111011111;
				8'b110001: c <= 9'b100000011;
				8'b1010111: c <= 9'b1010011;
				8'b1001110: c <= 9'b101110;
				8'b1101010: c <= 9'b101110001;
				8'b1001001: c <= 9'b100000010;
				8'b1100000: c <= 9'b1001111;
				8'b110111: c <= 9'b11001101;
				8'b1011101: c <= 9'b100011001;
				8'b1011011: c <= 9'b110000111;
				8'b111001: c <= 9'b10100;
				8'b1001010: c <= 9'b10100101;
				8'b110011: c <= 9'b10001001;
				8'b1101100: c <= 9'b11001111;
				8'b1110111: c <= 9'b1100111;
				8'b101011: c <= 9'b100000011;
				8'b1101011: c <= 9'b101101000;
				8'b111100: c <= 9'b100100101;
				8'b1000111: c <= 9'b1111001;
				8'b1011111: c <= 9'b11111011;
				8'b1110100: c <= 9'b1000100;
				8'b101101: c <= 9'b1001010;
				8'b1010011: c <= 9'b11111;
				8'b1100001: c <= 9'b11001000;
				8'b110101: c <= 9'b1000011;
				8'b1000100: c <= 9'b110001001;
				8'b1010001: c <= 9'b11101001;
				8'b1010100: c <= 9'b1100101;
				8'b1100110: c <= 9'b110100001;
				8'b101010: c <= 9'b111001111;
				8'b1011110: c <= 9'b111101111;
				8'b1100111: c <= 9'b11110101;
				8'b1011010: c <= 9'b111110011;
				8'b1000010: c <= 9'b111101;
				8'b111101: c <= 9'b110110100;
				8'b110000: c <= 9'b101100010;
				8'b111110: c <= 9'b110011;
				8'b1100010: c <= 9'b111011011;
				8'b1110000: c <= 9'b10111100;
				8'b1101001: c <= 9'b100000011;
				8'b1110011: c <= 9'b11110011;
				8'b1001100: c <= 9'b110010110;
				8'b100001: c <= 9'b100010000;
				8'b1000110: c <= 9'b1101010;
				8'b1110010: c <= 9'b111010100;
				8'b1010000: c <= 9'b10011000;
				8'b1111010: c <= 9'b10011011;
				8'b1010101: c <= 9'b111111010;
				8'b111011: c <= 9'b111011011;
				8'b1001101: c <= 9'b111100000;
				8'b111111: c <= 9'b11100010;
				8'b1101110: c <= 9'b10000;
				8'b1111011: c <= 9'b11001101;
				8'b1001011: c <= 9'b100011000;
				8'b1101111: c <= 9'b1001101;
				8'b1101000: c <= 9'b101;
				8'b101100: c <= 9'b110100011;
				8'b100100: c <= 9'b11111000;
				8'b1111000: c <= 9'b1001010;
				8'b1000101: c <= 9'b11110000;
				8'b1011001: c <= 9'b101101;
				8'b110100: c <= 9'b101110111;
				8'b1111001: c <= 9'b10100011;
				8'b1110001: c <= 9'b110001001;
				8'b1001111: c <= 9'b11000111;
				8'b1100101: c <= 9'b111111000;
				8'b1111110: c <= 9'b111010000;
				8'b1111100: c <= 9'b11110011;
				8'b1010110: c <= 9'b110001;
				8'b110010: c <= 9'b11100000;
				8'b1101101: c <= 9'b100111111;
				8'b100011: c <= 9'b111000100;
				8'b1110101: c <= 9'b1000000;
				8'b1111101: c <= 9'b100101011;
				8'b101001: c <= 9'b101101101;
				8'b1010010: c <= 9'b101010101;
				8'b1011000: c <= 9'b10110100;
				8'b101110: c <= 9'b1111101;
				8'b1000001: c <= 9'b101000100;
				default: c <= 9'b0;
			endcase
			9'b110011111 : case(di)
				8'b1000011: c <= 9'b1111011;
				8'b101000: c <= 9'b1010110;
				8'b111010: c <= 9'b10100110;
				8'b110110: c <= 9'b111010010;
				8'b1100100: c <= 9'b110001111;
				8'b1000000: c <= 9'b1101111;
				8'b1110110: c <= 9'b101;
				8'b100101: c <= 9'b101000110;
				8'b101111: c <= 9'b11111001;
				8'b100110: c <= 9'b10001001;
				8'b1100011: c <= 9'b1000011;
				8'b1001000: c <= 9'b101001001;
				8'b111000: c <= 9'b110101110;
				8'b110001: c <= 9'b101011101;
				8'b1010111: c <= 9'b100011111;
				8'b1001110: c <= 9'b110000111;
				8'b1101010: c <= 9'b100010100;
				8'b1001001: c <= 9'b10101101;
				8'b1100000: c <= 9'b11001001;
				8'b110111: c <= 9'b110101111;
				8'b1011101: c <= 9'b110010;
				8'b1011011: c <= 9'b10101101;
				8'b111001: c <= 9'b101010110;
				8'b1001010: c <= 9'b100001110;
				8'b110011: c <= 9'b101001001;
				8'b1101100: c <= 9'b101101001;
				8'b1110111: c <= 9'b1110001;
				8'b101011: c <= 9'b110111111;
				8'b1101011: c <= 9'b10000001;
				8'b111100: c <= 9'b11010111;
				8'b1000111: c <= 9'b100001101;
				8'b1011111: c <= 9'b110011100;
				8'b1110100: c <= 9'b1000001;
				8'b101101: c <= 9'b101110011;
				8'b1010011: c <= 9'b111100010;
				8'b1100001: c <= 9'b11101101;
				8'b110101: c <= 9'b1011001;
				8'b1000100: c <= 9'b10100011;
				8'b1010001: c <= 9'b11001010;
				8'b1010100: c <= 9'b10111101;
				8'b1100110: c <= 9'b11000011;
				8'b101010: c <= 9'b11000011;
				8'b1011110: c <= 9'b110000010;
				8'b1100111: c <= 9'b11000011;
				8'b1011010: c <= 9'b1;
				8'b1000010: c <= 9'b1000;
				8'b111101: c <= 9'b101101100;
				8'b110000: c <= 9'b100011111;
				8'b111110: c <= 9'b1101010;
				8'b1100010: c <= 9'b11010111;
				8'b1110000: c <= 9'b100110101;
				8'b1101001: c <= 9'b111100100;
				8'b1110011: c <= 9'b11010111;
				8'b1001100: c <= 9'b101111110;
				8'b100001: c <= 9'b110100100;
				8'b1000110: c <= 9'b10110001;
				8'b1110010: c <= 9'b10110111;
				8'b1010000: c <= 9'b101010001;
				8'b1111010: c <= 9'b10001000;
				8'b1010101: c <= 9'b101110110;
				8'b111011: c <= 9'b100100101;
				8'b1001101: c <= 9'b11110100;
				8'b111111: c <= 9'b100110010;
				8'b1101110: c <= 9'b111111101;
				8'b1111011: c <= 9'b100000101;
				8'b1001011: c <= 9'b1100;
				8'b1101111: c <= 9'b110001000;
				8'b1101000: c <= 9'b11001010;
				8'b101100: c <= 9'b1001000;
				8'b100100: c <= 9'b1001011;
				8'b1111000: c <= 9'b10010011;
				8'b1000101: c <= 9'b1101111;
				8'b1011001: c <= 9'b10011010;
				8'b110100: c <= 9'b101110001;
				8'b1111001: c <= 9'b101111110;
				8'b1110001: c <= 9'b1011;
				8'b1001111: c <= 9'b110111111;
				8'b1100101: c <= 9'b111010001;
				8'b1111110: c <= 9'b11011;
				8'b1111100: c <= 9'b110011100;
				8'b1010110: c <= 9'b100011011;
				8'b110010: c <= 9'b1100111;
				8'b1101101: c <= 9'b10111101;
				8'b100011: c <= 9'b11011000;
				8'b1110101: c <= 9'b10100011;
				8'b1111101: c <= 9'b101111000;
				8'b101001: c <= 9'b10010000;
				8'b1010010: c <= 9'b101011001;
				8'b1011000: c <= 9'b100101101;
				8'b101110: c <= 9'b10110010;
				8'b1000001: c <= 9'b10110001;
				default: c <= 9'b0;
			endcase
			9'b11111100 : case(di)
				8'b1000011: c <= 9'b100001011;
				8'b101000: c <= 9'b100100101;
				8'b111010: c <= 9'b10110011;
				8'b110110: c <= 9'b100000010;
				8'b1100100: c <= 9'b1111101;
				8'b1000000: c <= 9'b110100110;
				8'b1110110: c <= 9'b111100010;
				8'b100101: c <= 9'b110000011;
				8'b101111: c <= 9'b100100;
				8'b100110: c <= 9'b10000011;
				8'b1100011: c <= 9'b110011011;
				8'b1001000: c <= 9'b1101010;
				8'b111000: c <= 9'b111001;
				8'b110001: c <= 9'b11100;
				8'b1010111: c <= 9'b11001000;
				8'b1001110: c <= 9'b1010101;
				8'b1101010: c <= 9'b10001101;
				8'b1001001: c <= 9'b101011011;
				8'b1100000: c <= 9'b11100011;
				8'b110111: c <= 9'b1111110;
				8'b1011101: c <= 9'b111100110;
				8'b1011011: c <= 9'b101001001;
				8'b111001: c <= 9'b101011;
				8'b1001010: c <= 9'b1001000;
				8'b110011: c <= 9'b100101011;
				8'b1101100: c <= 9'b110010100;
				8'b1110111: c <= 9'b110111011;
				8'b101011: c <= 9'b110100111;
				8'b1101011: c <= 9'b101000110;
				8'b111100: c <= 9'b100000001;
				8'b1000111: c <= 9'b110101001;
				8'b1011111: c <= 9'b10010111;
				8'b1110100: c <= 9'b100111001;
				8'b101101: c <= 9'b11111011;
				8'b1010011: c <= 9'b101110000;
				8'b1100001: c <= 9'b11100111;
				8'b110101: c <= 9'b111000110;
				8'b1000100: c <= 9'b1000;
				8'b1010001: c <= 9'b11000000;
				8'b1010100: c <= 9'b111111111;
				8'b1100110: c <= 9'b101011101;
				8'b101010: c <= 9'b100101100;
				8'b1011110: c <= 9'b110100111;
				8'b1100111: c <= 9'b110110110;
				8'b1011010: c <= 9'b111111;
				8'b1000010: c <= 9'b100011010;
				8'b111101: c <= 9'b110100100;
				8'b110000: c <= 9'b11111110;
				8'b111110: c <= 9'b110100110;
				8'b1100010: c <= 9'b101101111;
				8'b1110000: c <= 9'b110010010;
				8'b1101001: c <= 9'b1011001;
				8'b1110011: c <= 9'b110010110;
				8'b1001100: c <= 9'b10101110;
				8'b100001: c <= 9'b10011001;
				8'b1000110: c <= 9'b11111110;
				8'b1110010: c <= 9'b10110101;
				8'b1010000: c <= 9'b110100100;
				8'b1111010: c <= 9'b110011001;
				8'b1010101: c <= 9'b11001010;
				8'b111011: c <= 9'b111011011;
				8'b1001101: c <= 9'b1000011;
				8'b111111: c <= 9'b101101010;
				8'b1101110: c <= 9'b111110011;
				8'b1111011: c <= 9'b11101001;
				8'b1001011: c <= 9'b10110011;
				8'b1101111: c <= 9'b10000011;
				8'b1101000: c <= 9'b1101;
				8'b101100: c <= 9'b101010101;
				8'b100100: c <= 9'b10110111;
				8'b1111000: c <= 9'b111000100;
				8'b1000101: c <= 9'b101100100;
				8'b1011001: c <= 9'b111;
				8'b110100: c <= 9'b10101111;
				8'b1111001: c <= 9'b11011100;
				8'b1110001: c <= 9'b101110000;
				8'b1001111: c <= 9'b1111011;
				8'b1100101: c <= 9'b1011;
				8'b1111110: c <= 9'b101110010;
				8'b1111100: c <= 9'b111000101;
				8'b1010110: c <= 9'b100110000;
				8'b110010: c <= 9'b11110111;
				8'b1101101: c <= 9'b111100100;
				8'b100011: c <= 9'b10100011;
				8'b1110101: c <= 9'b111110101;
				8'b1111101: c <= 9'b11111010;
				8'b101001: c <= 9'b11001100;
				8'b1010010: c <= 9'b110001000;
				8'b1011000: c <= 9'b101011111;
				8'b101110: c <= 9'b100110101;
				8'b1000001: c <= 9'b11110110;
				default: c <= 9'b0;
			endcase
			9'b100111010 : case(di)
				8'b1000011: c <= 9'b101101101;
				8'b101000: c <= 9'b11100100;
				8'b111010: c <= 9'b1111100;
				8'b110110: c <= 9'b111001101;
				8'b1100100: c <= 9'b101101101;
				8'b1000000: c <= 9'b10111101;
				8'b1110110: c <= 9'b10110101;
				8'b100101: c <= 9'b100101110;
				8'b101111: c <= 9'b1111100;
				8'b100110: c <= 9'b10010111;
				8'b1100011: c <= 9'b110101;
				8'b1001000: c <= 9'b1111110;
				8'b111000: c <= 9'b101101101;
				8'b110001: c <= 9'b101010100;
				8'b1010111: c <= 9'b101111001;
				8'b1001110: c <= 9'b1000001;
				8'b1101010: c <= 9'b11010;
				8'b1001001: c <= 9'b101100110;
				8'b1100000: c <= 9'b10001011;
				8'b110111: c <= 9'b101111001;
				8'b1011101: c <= 9'b100111101;
				8'b1011011: c <= 9'b111;
				8'b111001: c <= 9'b101010001;
				8'b1001010: c <= 9'b11100101;
				8'b110011: c <= 9'b100001011;
				8'b1101100: c <= 9'b11110101;
				8'b1110111: c <= 9'b110111110;
				8'b101011: c <= 9'b100100011;
				8'b1101011: c <= 9'b100010000;
				8'b111100: c <= 9'b11110110;
				8'b1000111: c <= 9'b110110101;
				8'b1011111: c <= 9'b11001101;
				8'b1110100: c <= 9'b100011;
				8'b101101: c <= 9'b10110111;
				8'b1010011: c <= 9'b100111100;
				8'b1100001: c <= 9'b100010;
				8'b110101: c <= 9'b111000011;
				8'b1000100: c <= 9'b1010010;
				8'b1010001: c <= 9'b1110101;
				8'b1010100: c <= 9'b111011;
				8'b1100110: c <= 9'b111010010;
				8'b101010: c <= 9'b110101111;
				8'b1011110: c <= 9'b1001001;
				8'b1100111: c <= 9'b111001101;
				8'b1011010: c <= 9'b1000100;
				8'b1000010: c <= 9'b1110001;
				8'b111101: c <= 9'b11100000;
				8'b110000: c <= 9'b111100011;
				8'b111110: c <= 9'b110101010;
				8'b1100010: c <= 9'b1011100;
				8'b1110000: c <= 9'b11111010;
				8'b1101001: c <= 9'b100010000;
				8'b1110011: c <= 9'b11010011;
				8'b1001100: c <= 9'b110001;
				8'b100001: c <= 9'b1110101;
				8'b1000110: c <= 9'b110101111;
				8'b1110010: c <= 9'b111010110;
				8'b1010000: c <= 9'b100011001;
				8'b1111010: c <= 9'b10111001;
				8'b1010101: c <= 9'b11000;
				8'b111011: c <= 9'b101011110;
				8'b1001101: c <= 9'b110100011;
				8'b111111: c <= 9'b100001001;
				8'b1101110: c <= 9'b1011000;
				8'b1111011: c <= 9'b11101011;
				8'b1001011: c <= 9'b1000111;
				8'b1101111: c <= 9'b101010111;
				8'b1101000: c <= 9'b10000101;
				8'b101100: c <= 9'b101101110;
				8'b100100: c <= 9'b10101100;
				8'b1111000: c <= 9'b101100101;
				8'b1000101: c <= 9'b100110;
				8'b1011001: c <= 9'b100100101;
				8'b110100: c <= 9'b110111100;
				8'b1111001: c <= 9'b100101101;
				8'b1110001: c <= 9'b10;
				8'b1001111: c <= 9'b10101110;
				8'b1100101: c <= 9'b11010000;
				8'b1111110: c <= 9'b1011;
				8'b1111100: c <= 9'b111010110;
				8'b1010110: c <= 9'b111110011;
				8'b110010: c <= 9'b101100110;
				8'b1101101: c <= 9'b1001;
				8'b100011: c <= 9'b10001101;
				8'b1110101: c <= 9'b1000110;
				8'b1111101: c <= 9'b10001001;
				8'b101001: c <= 9'b111011101;
				8'b1010010: c <= 9'b11000111;
				8'b1011000: c <= 9'b10000111;
				8'b101110: c <= 9'b101101;
				8'b1000001: c <= 9'b110101111;
				default: c <= 9'b0;
			endcase
			9'b101110001 : case(di)
				8'b1000011: c <= 9'b1110010;
				8'b101000: c <= 9'b101110110;
				8'b111010: c <= 9'b10101011;
				8'b110110: c <= 9'b1101001;
				8'b1100100: c <= 9'b1001110;
				8'b1000000: c <= 9'b111010;
				8'b1110110: c <= 9'b100011101;
				8'b100101: c <= 9'b100110111;
				8'b101111: c <= 9'b1100101;
				8'b100110: c <= 9'b111101100;
				8'b1100011: c <= 9'b110111010;
				8'b1001000: c <= 9'b110010001;
				8'b111000: c <= 9'b11110111;
				8'b110001: c <= 9'b11100001;
				8'b1010111: c <= 9'b101010100;
				8'b1001110: c <= 9'b100100011;
				8'b1101010: c <= 9'b110001000;
				8'b1001001: c <= 9'b100010100;
				8'b1100000: c <= 9'b10111100;
				8'b110111: c <= 9'b101101110;
				8'b1011101: c <= 9'b1100;
				8'b1011011: c <= 9'b101101011;
				8'b111001: c <= 9'b11001000;
				8'b1001010: c <= 9'b110001101;
				8'b110011: c <= 9'b110110111;
				8'b1101100: c <= 9'b111101000;
				8'b1110111: c <= 9'b100111000;
				8'b101011: c <= 9'b10100101;
				8'b1101011: c <= 9'b101110111;
				8'b111100: c <= 9'b100010110;
				8'b1000111: c <= 9'b101111110;
				8'b1011111: c <= 9'b111111110;
				8'b1110100: c <= 9'b1010010;
				8'b101101: c <= 9'b111111000;
				8'b1010011: c <= 9'b1001000;
				8'b1100001: c <= 9'b110100110;
				8'b110101: c <= 9'b110000;
				8'b1000100: c <= 9'b101100001;
				8'b1010001: c <= 9'b101000100;
				8'b1010100: c <= 9'b11010111;
				8'b1100110: c <= 9'b111111;
				8'b101010: c <= 9'b100000001;
				8'b1011110: c <= 9'b110110100;
				8'b1100111: c <= 9'b100110;
				8'b1011010: c <= 9'b10001010;
				8'b1000010: c <= 9'b10101000;
				8'b111101: c <= 9'b111010000;
				8'b110000: c <= 9'b101110001;
				8'b111110: c <= 9'b110110;
				8'b1100010: c <= 9'b10111110;
				8'b1110000: c <= 9'b11011000;
				8'b1101001: c <= 9'b100000101;
				8'b1110011: c <= 9'b1111111;
				8'b1001100: c <= 9'b111011011;
				8'b100001: c <= 9'b1110100;
				8'b1000110: c <= 9'b11111010;
				8'b1110010: c <= 9'b101101000;
				8'b1010000: c <= 9'b100100110;
				8'b1111010: c <= 9'b11111000;
				8'b1010101: c <= 9'b111011101;
				8'b111011: c <= 9'b1011011;
				8'b1001101: c <= 9'b11110100;
				8'b111111: c <= 9'b101000111;
				8'b1101110: c <= 9'b110011110;
				8'b1111011: c <= 9'b1001000;
				8'b1001011: c <= 9'b11011;
				8'b1101111: c <= 9'b111110110;
				8'b1101000: c <= 9'b10001001;
				8'b101100: c <= 9'b1011;
				8'b100100: c <= 9'b1000101;
				8'b1111000: c <= 9'b101010010;
				8'b1000101: c <= 9'b111011110;
				8'b1011001: c <= 9'b1100010;
				8'b110100: c <= 9'b1100001;
				8'b1111001: c <= 9'b110001000;
				8'b1110001: c <= 9'b10001101;
				8'b1001111: c <= 9'b10101010;
				8'b1100101: c <= 9'b111100001;
				8'b1111110: c <= 9'b11111001;
				8'b1111100: c <= 9'b110110110;
				8'b1010110: c <= 9'b1010001;
				8'b110010: c <= 9'b10000010;
				8'b1101101: c <= 9'b11000000;
				8'b100011: c <= 9'b100100111;
				8'b1110101: c <= 9'b1101111;
				8'b1111101: c <= 9'b10100011;
				8'b101001: c <= 9'b111001111;
				8'b1010010: c <= 9'b110110101;
				8'b1011000: c <= 9'b111001;
				8'b101110: c <= 9'b100101;
				8'b1000001: c <= 9'b101010110;
				default: c <= 9'b0;
			endcase
			9'b110110 : case(di)
				8'b1000011: c <= 9'b111111110;
				8'b101000: c <= 9'b11100101;
				8'b111010: c <= 9'b100010101;
				8'b110110: c <= 9'b1101001;
				8'b1100100: c <= 9'b100000100;
				8'b1000000: c <= 9'b110011110;
				8'b1110110: c <= 9'b100110111;
				8'b100101: c <= 9'b101001110;
				8'b101111: c <= 9'b11010010;
				8'b100110: c <= 9'b10001001;
				8'b1100011: c <= 9'b101110111;
				8'b1001000: c <= 9'b100000001;
				8'b111000: c <= 9'b111010010;
				8'b110001: c <= 9'b110100010;
				8'b1010111: c <= 9'b101110000;
				8'b1001110: c <= 9'b100100110;
				8'b1101010: c <= 9'b101111000;
				8'b1001001: c <= 9'b100010010;
				8'b1100000: c <= 9'b101100100;
				8'b110111: c <= 9'b111100;
				8'b1011101: c <= 9'b10101111;
				8'b1011011: c <= 9'b1001011;
				8'b111001: c <= 9'b111101010;
				8'b1001010: c <= 9'b10110010;
				8'b110011: c <= 9'b1111010;
				8'b1101100: c <= 9'b110100001;
				8'b1110111: c <= 9'b1000111;
				8'b101011: c <= 9'b1110011;
				8'b1101011: c <= 9'b11111;
				8'b111100: c <= 9'b101111000;
				8'b1000111: c <= 9'b100111110;
				8'b1011111: c <= 9'b10110111;
				8'b1110100: c <= 9'b110101101;
				8'b101101: c <= 9'b110001001;
				8'b1010011: c <= 9'b10110101;
				8'b1100001: c <= 9'b111011010;
				8'b110101: c <= 9'b110111100;
				8'b1000100: c <= 9'b100011;
				8'b1010001: c <= 9'b10010111;
				8'b1010100: c <= 9'b11011001;
				8'b1100110: c <= 9'b1111010;
				8'b101010: c <= 9'b1100100;
				8'b1011110: c <= 9'b1011100;
				8'b1100111: c <= 9'b110001000;
				8'b1011010: c <= 9'b10011011;
				8'b1000010: c <= 9'b111110011;
				8'b111101: c <= 9'b100011011;
				8'b110000: c <= 9'b11100011;
				8'b111110: c <= 9'b110011011;
				8'b1100010: c <= 9'b1000100;
				8'b1110000: c <= 9'b100110101;
				8'b1101001: c <= 9'b1101000;
				8'b1110011: c <= 9'b1000100;
				8'b1001100: c <= 9'b11011001;
				8'b100001: c <= 9'b11110110;
				8'b1000110: c <= 9'b111110101;
				8'b1110010: c <= 9'b10111010;
				8'b1010000: c <= 9'b101011011;
				8'b1111010: c <= 9'b100001010;
				8'b1010101: c <= 9'b1100110;
				8'b111011: c <= 9'b111;
				8'b1001101: c <= 9'b100001011;
				8'b111111: c <= 9'b101101010;
				8'b1101110: c <= 9'b110110110;
				8'b1111011: c <= 9'b100001111;
				8'b1001011: c <= 9'b101001100;
				8'b1101111: c <= 9'b1000010;
				8'b1101000: c <= 9'b110111011;
				8'b101100: c <= 9'b111000100;
				8'b100100: c <= 9'b111100101;
				8'b1111000: c <= 9'b111011100;
				8'b1000101: c <= 9'b111110001;
				8'b1011001: c <= 9'b10101011;
				8'b110100: c <= 9'b10111011;
				8'b1111001: c <= 9'b11000011;
				8'b1110001: c <= 9'b1100100;
				8'b1001111: c <= 9'b100010100;
				8'b1100101: c <= 9'b10101011;
				8'b1111110: c <= 9'b111000011;
				8'b1111100: c <= 9'b110000101;
				8'b1010110: c <= 9'b101010010;
				8'b110010: c <= 9'b10110110;
				8'b1101101: c <= 9'b1100100;
				8'b100011: c <= 9'b1111;
				8'b1110101: c <= 9'b11000110;
				8'b1111101: c <= 9'b10010111;
				8'b101001: c <= 9'b110001001;
				8'b1010010: c <= 9'b111101101;
				8'b1011000: c <= 9'b100111;
				8'b101110: c <= 9'b101010;
				8'b1000001: c <= 9'b111000000;
				default: c <= 9'b0;
			endcase
			9'b11100011 : case(di)
				8'b1000011: c <= 9'b110100001;
				8'b101000: c <= 9'b100110101;
				8'b111010: c <= 9'b1;
				8'b110110: c <= 9'b101100000;
				8'b1100100: c <= 9'b101110;
				8'b1000000: c <= 9'b1010001;
				8'b1110110: c <= 9'b110000011;
				8'b100101: c <= 9'b1010000;
				8'b101111: c <= 9'b111000101;
				8'b100110: c <= 9'b110011001;
				8'b1100011: c <= 9'b100111101;
				8'b1001000: c <= 9'b111001001;
				8'b111000: c <= 9'b111001000;
				8'b110001: c <= 9'b10010100;
				8'b1010111: c <= 9'b10110100;
				8'b1001110: c <= 9'b111001010;
				8'b1101010: c <= 9'b111000111;
				8'b1001001: c <= 9'b101101;
				8'b1100000: c <= 9'b111110001;
				8'b110111: c <= 9'b11000;
				8'b1011101: c <= 9'b1001110;
				8'b1011011: c <= 9'b11010100;
				8'b111001: c <= 9'b11001101;
				8'b1001010: c <= 9'b10011101;
				8'b110011: c <= 9'b1111;
				8'b1101100: c <= 9'b1000011;
				8'b1110111: c <= 9'b110011011;
				8'b101011: c <= 9'b110001110;
				8'b1101011: c <= 9'b101110111;
				8'b111100: c <= 9'b111010100;
				8'b1000111: c <= 9'b1110;
				8'b1011111: c <= 9'b11001000;
				8'b1110100: c <= 9'b10010111;
				8'b101101: c <= 9'b111100010;
				8'b1010011: c <= 9'b11101000;
				8'b1100001: c <= 9'b11010001;
				8'b110101: c <= 9'b11111011;
				8'b1000100: c <= 9'b111100010;
				8'b1010001: c <= 9'b111101111;
				8'b1010100: c <= 9'b10000011;
				8'b1100110: c <= 9'b101000100;
				8'b101010: c <= 9'b101101100;
				8'b1011110: c <= 9'b1100101;
				8'b1100111: c <= 9'b111100010;
				8'b1011010: c <= 9'b10001011;
				8'b1000010: c <= 9'b110111110;
				8'b111101: c <= 9'b111101110;
				8'b110000: c <= 9'b111101111;
				8'b111110: c <= 9'b101100110;
				8'b1100010: c <= 9'b1111000;
				8'b1110000: c <= 9'b100101100;
				8'b1101001: c <= 9'b100110011;
				8'b1110011: c <= 9'b111111011;
				8'b1001100: c <= 9'b111010001;
				8'b100001: c <= 9'b10101011;
				8'b1000110: c <= 9'b111101101;
				8'b1110010: c <= 9'b111111;
				8'b1010000: c <= 9'b10001000;
				8'b1111010: c <= 9'b111000111;
				8'b1010101: c <= 9'b10011010;
				8'b111011: c <= 9'b100111111;
				8'b1001101: c <= 9'b11010;
				8'b111111: c <= 9'b100010000;
				8'b1101110: c <= 9'b101010100;
				8'b1111011: c <= 9'b10110;
				8'b1001011: c <= 9'b101011110;
				8'b1101111: c <= 9'b101001001;
				8'b1101000: c <= 9'b1011100;
				8'b101100: c <= 9'b11100;
				8'b100100: c <= 9'b111010111;
				8'b1111000: c <= 9'b100111011;
				8'b1000101: c <= 9'b10111110;
				8'b1011001: c <= 9'b111000000;
				8'b110100: c <= 9'b100011000;
				8'b1111001: c <= 9'b1000111;
				8'b1110001: c <= 9'b101010010;
				8'b1001111: c <= 9'b101111001;
				8'b1100101: c <= 9'b110000110;
				8'b1111110: c <= 9'b110010011;
				8'b1111100: c <= 9'b110010;
				8'b1010110: c <= 9'b110101;
				8'b110010: c <= 9'b11010001;
				8'b1101101: c <= 9'b1011010;
				8'b100011: c <= 9'b111111101;
				8'b1110101: c <= 9'b1010010;
				8'b1111101: c <= 9'b110100011;
				8'b101001: c <= 9'b10001111;
				8'b1010010: c <= 9'b111000000;
				8'b1011000: c <= 9'b111111000;
				8'b101110: c <= 9'b110000110;
				8'b1000001: c <= 9'b111011;
				default: c <= 9'b0;
			endcase
			9'b110101 : case(di)
				8'b1000011: c <= 9'b110011101;
				8'b101000: c <= 9'b101011;
				8'b111010: c <= 9'b100111101;
				8'b110110: c <= 9'b100010110;
				8'b1100100: c <= 9'b10111111;
				8'b1000000: c <= 9'b10011010;
				8'b1110110: c <= 9'b111001001;
				8'b100101: c <= 9'b11101000;
				8'b101111: c <= 9'b1110001;
				8'b100110: c <= 9'b1101111;
				8'b1100011: c <= 9'b1000001;
				8'b1001000: c <= 9'b111010111;
				8'b111000: c <= 9'b101101;
				8'b110001: c <= 9'b100111111;
				8'b1010111: c <= 9'b1100111;
				8'b1001110: c <= 9'b101110;
				8'b1101010: c <= 9'b100000001;
				8'b1001001: c <= 9'b1100001;
				8'b1100000: c <= 9'b100010000;
				8'b110111: c <= 9'b110001100;
				8'b1011101: c <= 9'b10000111;
				8'b1011011: c <= 9'b110101100;
				8'b111001: c <= 9'b111101101;
				8'b1001010: c <= 9'b110111111;
				8'b110011: c <= 9'b101110000;
				8'b1101100: c <= 9'b101010011;
				8'b1110111: c <= 9'b101001011;
				8'b101011: c <= 9'b10011100;
				8'b1101011: c <= 9'b10101111;
				8'b111100: c <= 9'b101101011;
				8'b1000111: c <= 9'b11001110;
				8'b1011111: c <= 9'b11110100;
				8'b1110100: c <= 9'b110101001;
				8'b101101: c <= 9'b111011111;
				8'b1010011: c <= 9'b100010110;
				8'b1100001: c <= 9'b11011011;
				8'b110101: c <= 9'b10010101;
				8'b1000100: c <= 9'b1011001;
				8'b1010001: c <= 9'b10100011;
				8'b1010100: c <= 9'b11100100;
				8'b1100110: c <= 9'b11111101;
				8'b101010: c <= 9'b1110010;
				8'b1011110: c <= 9'b101011000;
				8'b1100111: c <= 9'b110100;
				8'b1011010: c <= 9'b111110001;
				8'b1000010: c <= 9'b11110101;
				8'b111101: c <= 9'b11100100;
				8'b110000: c <= 9'b110100110;
				8'b111110: c <= 9'b111000100;
				8'b1100010: c <= 9'b1000101;
				8'b1110000: c <= 9'b101001110;
				8'b1101001: c <= 9'b10101110;
				8'b1110011: c <= 9'b11111001;
				8'b1001100: c <= 9'b11111000;
				8'b100001: c <= 9'b11111;
				8'b1000110: c <= 9'b11110111;
				8'b1110010: c <= 9'b11001101;
				8'b1010000: c <= 9'b101111110;
				8'b1111010: c <= 9'b10011010;
				8'b1010101: c <= 9'b101110011;
				8'b111011: c <= 9'b100101110;
				8'b1001101: c <= 9'b1111110;
				8'b111111: c <= 9'b1001;
				8'b1101110: c <= 9'b111001010;
				8'b1111011: c <= 9'b100001011;
				8'b1001011: c <= 9'b11010100;
				8'b1101111: c <= 9'b1100111;
				8'b1101000: c <= 9'b100010101;
				8'b101100: c <= 9'b100000101;
				8'b100100: c <= 9'b101101101;
				8'b1111000: c <= 9'b10001011;
				8'b1000101: c <= 9'b101000110;
				8'b1011001: c <= 9'b11100010;
				8'b110100: c <= 9'b110110010;
				8'b1111001: c <= 9'b11111011;
				8'b1110001: c <= 9'b1011110;
				8'b1001111: c <= 9'b111;
				8'b1100101: c <= 9'b10101111;
				8'b1111110: c <= 9'b1101001;
				8'b1111100: c <= 9'b110011111;
				8'b1010110: c <= 9'b111000101;
				8'b110010: c <= 9'b101110000;
				8'b1101101: c <= 9'b10001011;
				8'b100011: c <= 9'b1111000;
				8'b1110101: c <= 9'b100001111;
				8'b1111101: c <= 9'b110010101;
				8'b101001: c <= 9'b10110001;
				8'b1010010: c <= 9'b101010011;
				8'b1011000: c <= 9'b101101010;
				8'b101110: c <= 9'b100111111;
				8'b1000001: c <= 9'b1101110;
				default: c <= 9'b0;
			endcase
			9'b101111000 : case(di)
				8'b1000011: c <= 9'b110101011;
				8'b101000: c <= 9'b110111110;
				8'b111010: c <= 9'b10111110;
				8'b110110: c <= 9'b1110011;
				8'b1100100: c <= 9'b10000101;
				8'b1000000: c <= 9'b110101010;
				8'b1110110: c <= 9'b10110111;
				8'b100101: c <= 9'b110001001;
				8'b101111: c <= 9'b111101101;
				8'b100110: c <= 9'b10011010;
				8'b1100011: c <= 9'b101011101;
				8'b1001000: c <= 9'b11101101;
				8'b111000: c <= 9'b11000110;
				8'b110001: c <= 9'b1111101;
				8'b1010111: c <= 9'b101100110;
				8'b1001110: c <= 9'b10110111;
				8'b1101010: c <= 9'b100000100;
				8'b1001001: c <= 9'b110000001;
				8'b1100000: c <= 9'b1011100;
				8'b110111: c <= 9'b101111111;
				8'b1011101: c <= 9'b10001110;
				8'b1011011: c <= 9'b101111001;
				8'b111001: c <= 9'b11011101;
				8'b1001010: c <= 9'b1001110;
				8'b110011: c <= 9'b101011101;
				8'b1101100: c <= 9'b10110;
				8'b1110111: c <= 9'b10011001;
				8'b101011: c <= 9'b111;
				8'b1101011: c <= 9'b1000;
				8'b111100: c <= 9'b10110010;
				8'b1000111: c <= 9'b10010011;
				8'b1011111: c <= 9'b10111010;
				8'b1110100: c <= 9'b101101111;
				8'b101101: c <= 9'b101010010;
				8'b1010011: c <= 9'b10000110;
				8'b1100001: c <= 9'b111110011;
				8'b110101: c <= 9'b100111011;
				8'b1000100: c <= 9'b1010011;
				8'b1010001: c <= 9'b110001111;
				8'b1010100: c <= 9'b111011001;
				8'b1100110: c <= 9'b11011011;
				8'b101010: c <= 9'b10111100;
				8'b1011110: c <= 9'b110100011;
				8'b1100111: c <= 9'b11100111;
				8'b1011010: c <= 9'b10100011;
				8'b1000010: c <= 9'b101000110;
				8'b111101: c <= 9'b11011000;
				8'b110000: c <= 9'b110000110;
				8'b111110: c <= 9'b1011111;
				8'b1100010: c <= 9'b110110000;
				8'b1110000: c <= 9'b11010001;
				8'b1101001: c <= 9'b110100111;
				8'b1110011: c <= 9'b111111101;
				8'b1001100: c <= 9'b111111001;
				8'b100001: c <= 9'b100110100;
				8'b1000110: c <= 9'b110010100;
				8'b1110010: c <= 9'b110011011;
				8'b1010000: c <= 9'b111000100;
				8'b1111010: c <= 9'b100101011;
				8'b1010101: c <= 9'b1100111;
				8'b111011: c <= 9'b101100;
				8'b1001101: c <= 9'b1101;
				8'b111111: c <= 9'b101;
				8'b1101110: c <= 9'b11010001;
				8'b1111011: c <= 9'b111101000;
				8'b1001011: c <= 9'b111010110;
				8'b1101111: c <= 9'b11111000;
				8'b1101000: c <= 9'b11011010;
				8'b101100: c <= 9'b11110110;
				8'b100100: c <= 9'b10101001;
				8'b1111000: c <= 9'b100111000;
				8'b1000101: c <= 9'b110101010;
				8'b1011001: c <= 9'b110000110;
				8'b110100: c <= 9'b100000001;
				8'b1111001: c <= 9'b11110;
				8'b1110001: c <= 9'b1100010;
				8'b1001111: c <= 9'b1000100;
				8'b1100101: c <= 9'b100011010;
				8'b1111110: c <= 9'b111001;
				8'b1111100: c <= 9'b100101000;
				8'b1010110: c <= 9'b11100101;
				8'b110010: c <= 9'b100100;
				8'b1101101: c <= 9'b100100;
				8'b100011: c <= 9'b100100101;
				8'b1110101: c <= 9'b110110011;
				8'b1111101: c <= 9'b1110001;
				8'b101001: c <= 9'b10100110;
				8'b1010010: c <= 9'b10110110;
				8'b1011000: c <= 9'b100111;
				8'b101110: c <= 9'b101110011;
				8'b1000001: c <= 9'b100000101;
				default: c <= 9'b0;
			endcase
			9'b100 : case(di)
				8'b1000011: c <= 9'b10101101;
				8'b101000: c <= 9'b111010100;
				8'b111010: c <= 9'b10111001;
				8'b110110: c <= 9'b101001111;
				8'b1100100: c <= 9'b101010111;
				8'b1000000: c <= 9'b11000110;
				8'b1110110: c <= 9'b110111;
				8'b100101: c <= 9'b100101;
				8'b101111: c <= 9'b100000010;
				8'b100110: c <= 9'b100011000;
				8'b1100011: c <= 9'b10000110;
				8'b1001000: c <= 9'b11100;
				8'b111000: c <= 9'b1010001;
				8'b110001: c <= 9'b1000010;
				8'b1010111: c <= 9'b101010010;
				8'b1001110: c <= 9'b11011;
				8'b1101010: c <= 9'b100010100;
				8'b1001001: c <= 9'b10000010;
				8'b1100000: c <= 9'b101100000;
				8'b110111: c <= 9'b101010100;
				8'b1011101: c <= 9'b10001110;
				8'b1011011: c <= 9'b10010101;
				8'b111001: c <= 9'b1100110;
				8'b1001010: c <= 9'b110010010;
				8'b110011: c <= 9'b111111111;
				8'b1101100: c <= 9'b110101101;
				8'b1110111: c <= 9'b111000100;
				8'b101011: c <= 9'b10110001;
				8'b1101011: c <= 9'b11110111;
				8'b111100: c <= 9'b11101001;
				8'b1000111: c <= 9'b1000000;
				8'b1011111: c <= 9'b111011;
				8'b1110100: c <= 9'b11111000;
				8'b101101: c <= 9'b110011010;
				8'b1010011: c <= 9'b100001111;
				8'b1100001: c <= 9'b110011110;
				8'b110101: c <= 9'b110110000;
				8'b1000100: c <= 9'b110001011;
				8'b1010001: c <= 9'b100111010;
				8'b1010100: c <= 9'b11001000;
				8'b1100110: c <= 9'b1000010;
				8'b101010: c <= 9'b10101111;
				8'b1011110: c <= 9'b100001111;
				8'b1100111: c <= 9'b101001011;
				8'b1011010: c <= 9'b111101000;
				8'b1000010: c <= 9'b101110101;
				8'b111101: c <= 9'b10111101;
				8'b110000: c <= 9'b110100001;
				8'b111110: c <= 9'b110;
				8'b1100010: c <= 9'b11111000;
				8'b1110000: c <= 9'b1111010;
				8'b1101001: c <= 9'b1110011;
				8'b1110011: c <= 9'b111011101;
				8'b1001100: c <= 9'b101111111;
				8'b100001: c <= 9'b101000111;
				8'b1000110: c <= 9'b110111011;
				8'b1110010: c <= 9'b1000000;
				8'b1010000: c <= 9'b100110011;
				8'b1111010: c <= 9'b100101011;
				8'b1010101: c <= 9'b10100011;
				8'b111011: c <= 9'b111010100;
				8'b1001101: c <= 9'b10101011;
				8'b111111: c <= 9'b10111000;
				8'b1101110: c <= 9'b11001001;
				8'b1111011: c <= 9'b10000010;
				8'b1001011: c <= 9'b101110100;
				8'b1101111: c <= 9'b1111001;
				8'b1101000: c <= 9'b11110010;
				8'b101100: c <= 9'b101100010;
				8'b100100: c <= 9'b101110010;
				8'b1111000: c <= 9'b111111101;
				8'b1000101: c <= 9'b10000;
				8'b1011001: c <= 9'b11010101;
				8'b110100: c <= 9'b110011001;
				8'b1111001: c <= 9'b101111111;
				8'b1110001: c <= 9'b11010111;
				8'b1001111: c <= 9'b110100001;
				8'b1100101: c <= 9'b111101;
				8'b1111110: c <= 9'b111000011;
				8'b1111100: c <= 9'b100010001;
				8'b1010110: c <= 9'b111111110;
				8'b110010: c <= 9'b10010001;
				8'b1101101: c <= 9'b111101001;
				8'b100011: c <= 9'b1111110;
				8'b1110101: c <= 9'b10111011;
				8'b1111101: c <= 9'b111111101;
				8'b101001: c <= 9'b110001000;
				8'b1010010: c <= 9'b11111000;
				8'b1011000: c <= 9'b110000111;
				8'b101110: c <= 9'b1011;
				8'b1000001: c <= 9'b111111111;
				default: c <= 9'b0;
			endcase
			9'b110001110 : case(di)
				8'b1000011: c <= 9'b10011011;
				8'b101000: c <= 9'b111111011;
				8'b111010: c <= 9'b101110;
				8'b110110: c <= 9'b1010110;
				8'b1100100: c <= 9'b100100000;
				8'b1000000: c <= 9'b100010001;
				8'b1110110: c <= 9'b10010101;
				8'b100101: c <= 9'b111111;
				8'b101111: c <= 9'b111011110;
				8'b100110: c <= 9'b100101101;
				8'b1100011: c <= 9'b101100000;
				8'b1001000: c <= 9'b101110000;
				8'b111000: c <= 9'b100101011;
				8'b110001: c <= 9'b11010001;
				8'b1010111: c <= 9'b1000110;
				8'b1001110: c <= 9'b110110101;
				8'b1101010: c <= 9'b10000000;
				8'b1001001: c <= 9'b10101101;
				8'b1100000: c <= 9'b110000;
				8'b110111: c <= 9'b111100000;
				8'b1011101: c <= 9'b110010111;
				8'b1011011: c <= 9'b10110101;
				8'b111001: c <= 9'b100;
				8'b1001010: c <= 9'b1111;
				8'b110011: c <= 9'b10000;
				8'b1101100: c <= 9'b1010111;
				8'b1110111: c <= 9'b11010011;
				8'b101011: c <= 9'b101010101;
				8'b1101011: c <= 9'b10010111;
				8'b111100: c <= 9'b10110;
				8'b1000111: c <= 9'b1110001;
				8'b1011111: c <= 9'b1000101;
				8'b1110100: c <= 9'b100100;
				8'b101101: c <= 9'b100001100;
				8'b1010011: c <= 9'b10101001;
				8'b1100001: c <= 9'b111100011;
				8'b110101: c <= 9'b100111;
				8'b1000100: c <= 9'b11011010;
				8'b1010001: c <= 9'b1001100;
				8'b1010100: c <= 9'b1011010;
				8'b1100110: c <= 9'b111011;
				8'b101010: c <= 9'b110011111;
				8'b1011110: c <= 9'b110000110;
				8'b1100111: c <= 9'b111011011;
				8'b1011010: c <= 9'b11110011;
				8'b1000010: c <= 9'b100100111;
				8'b111101: c <= 9'b10001010;
				8'b110000: c <= 9'b11110111;
				8'b111110: c <= 9'b101001010;
				8'b1100010: c <= 9'b110001011;
				8'b1110000: c <= 9'b100011100;
				8'b1101001: c <= 9'b1011011;
				8'b1110011: c <= 9'b101110100;
				8'b1001100: c <= 9'b100100;
				8'b100001: c <= 9'b110001011;
				8'b1000110: c <= 9'b100111111;
				8'b1110010: c <= 9'b11000111;
				8'b1010000: c <= 9'b110100111;
				8'b1111010: c <= 9'b11111100;
				8'b1010101: c <= 9'b111001010;
				8'b111011: c <= 9'b111000010;
				8'b1001101: c <= 9'b101100100;
				8'b111111: c <= 9'b110111010;
				8'b1101110: c <= 9'b1010001;
				8'b1111011: c <= 9'b10001010;
				8'b1001011: c <= 9'b111001101;
				8'b1101111: c <= 9'b110101101;
				8'b1101000: c <= 9'b111100011;
				8'b101100: c <= 9'b10111111;
				8'b100100: c <= 9'b10000000;
				8'b1111000: c <= 9'b110000110;
				8'b1000101: c <= 9'b10010111;
				8'b1011001: c <= 9'b101001;
				8'b110100: c <= 9'b100110010;
				8'b1111001: c <= 9'b100011101;
				8'b1110001: c <= 9'b100;
				8'b1001111: c <= 9'b101011111;
				8'b1100101: c <= 9'b1110101;
				8'b1111110: c <= 9'b100110;
				8'b1111100: c <= 9'b110110000;
				8'b1010110: c <= 9'b10100110;
				8'b110010: c <= 9'b111011111;
				8'b1101101: c <= 9'b101100000;
				8'b100011: c <= 9'b111011010;
				8'b1110101: c <= 9'b101000;
				8'b1111101: c <= 9'b10100011;
				8'b101001: c <= 9'b111100010;
				8'b1010010: c <= 9'b1;
				8'b1011000: c <= 9'b10111000;
				8'b101110: c <= 9'b10111101;
				8'b1000001: c <= 9'b10010100;
				default: c <= 9'b0;
			endcase
			9'b11110010 : case(di)
				8'b1000011: c <= 9'b11011;
				8'b101000: c <= 9'b100011111;
				8'b111010: c <= 9'b101001001;
				8'b110110: c <= 9'b101000011;
				8'b1100100: c <= 9'b1100101;
				8'b1000000: c <= 9'b1000010;
				8'b1110110: c <= 9'b11110;
				8'b100101: c <= 9'b1001;
				8'b101111: c <= 9'b111101100;
				8'b100110: c <= 9'b10110010;
				8'b1100011: c <= 9'b101000011;
				8'b1001000: c <= 9'b100111011;
				8'b111000: c <= 9'b111001100;
				8'b110001: c <= 9'b11010000;
				8'b1010111: c <= 9'b101110;
				8'b1001110: c <= 9'b100001;
				8'b1101010: c <= 9'b100111010;
				8'b1001001: c <= 9'b10011101;
				8'b1100000: c <= 9'b11110010;
				8'b110111: c <= 9'b111011100;
				8'b1011101: c <= 9'b10011;
				8'b1011011: c <= 9'b101010011;
				8'b111001: c <= 9'b110001101;
				8'b1001010: c <= 9'b11010100;
				8'b110011: c <= 9'b111101111;
				8'b1101100: c <= 9'b10100011;
				8'b1110111: c <= 9'b1101000;
				8'b101011: c <= 9'b10000010;
				8'b1101011: c <= 9'b111011;
				8'b111100: c <= 9'b111110011;
				8'b1000111: c <= 9'b100100111;
				8'b1011111: c <= 9'b100011;
				8'b1110100: c <= 9'b100110011;
				8'b101101: c <= 9'b1101110;
				8'b1010011: c <= 9'b101000001;
				8'b1100001: c <= 9'b1100111;
				8'b110101: c <= 9'b1100100;
				8'b1000100: c <= 9'b101001100;
				8'b1010001: c <= 9'b1001111;
				8'b1010100: c <= 9'b111010111;
				8'b1100110: c <= 9'b10010000;
				8'b101010: c <= 9'b11110;
				8'b1011110: c <= 9'b111110110;
				8'b1100111: c <= 9'b1001111;
				8'b1011010: c <= 9'b11000011;
				8'b1000010: c <= 9'b110111000;
				8'b111101: c <= 9'b100110111;
				8'b110000: c <= 9'b111101101;
				8'b111110: c <= 9'b100011001;
				8'b1100010: c <= 9'b101010100;
				8'b1110000: c <= 9'b11100011;
				8'b1101001: c <= 9'b11000110;
				8'b1110011: c <= 9'b110010101;
				8'b1001100: c <= 9'b100101000;
				8'b100001: c <= 9'b11111110;
				8'b1000110: c <= 9'b110111010;
				8'b1110010: c <= 9'b110100000;
				8'b1010000: c <= 9'b101110100;
				8'b1111010: c <= 9'b11110011;
				8'b1010101: c <= 9'b11000100;
				8'b111011: c <= 9'b101110101;
				8'b1001101: c <= 9'b10010001;
				8'b111111: c <= 9'b1110001;
				8'b1101110: c <= 9'b101101110;
				8'b1111011: c <= 9'b110010010;
				8'b1001011: c <= 9'b101;
				8'b1101111: c <= 9'b100100000;
				8'b1101000: c <= 9'b101001111;
				8'b101100: c <= 9'b100111000;
				8'b100100: c <= 9'b101110101;
				8'b1111000: c <= 9'b110101;
				8'b1000101: c <= 9'b10001111;
				8'b1011001: c <= 9'b1011001;
				8'b110100: c <= 9'b101010001;
				8'b1111001: c <= 9'b101010111;
				8'b1110001: c <= 9'b100011010;
				8'b1001111: c <= 9'b111011010;
				8'b1100101: c <= 9'b101000;
				8'b1111110: c <= 9'b10111000;
				8'b1111100: c <= 9'b10001011;
				8'b1010110: c <= 9'b110001111;
				8'b110010: c <= 9'b110010101;
				8'b1101101: c <= 9'b1000011;
				8'b100011: c <= 9'b11101111;
				8'b1110101: c <= 9'b11110000;
				8'b1111101: c <= 9'b100000110;
				8'b101001: c <= 9'b1001;
				8'b1010010: c <= 9'b10010001;
				8'b1011000: c <= 9'b10010000;
				8'b101110: c <= 9'b101101100;
				8'b1000001: c <= 9'b111010;
				default: c <= 9'b0;
			endcase
			9'b110010110 : case(di)
				8'b1000011: c <= 9'b1100111;
				8'b101000: c <= 9'b111111;
				8'b111010: c <= 9'b1000110;
				8'b110110: c <= 9'b101000;
				8'b1100100: c <= 9'b100111011;
				8'b1000000: c <= 9'b10101;
				8'b1110110: c <= 9'b10110110;
				8'b100101: c <= 9'b110101111;
				8'b101111: c <= 9'b100;
				8'b100110: c <= 9'b111100110;
				8'b1100011: c <= 9'b100110111;
				8'b1001000: c <= 9'b101010011;
				8'b111000: c <= 9'b11100110;
				8'b110001: c <= 9'b101101001;
				8'b1010111: c <= 9'b11100101;
				8'b1001110: c <= 9'b110011000;
				8'b1101010: c <= 9'b1111011;
				8'b1001001: c <= 9'b11001001;
				8'b1100000: c <= 9'b101101100;
				8'b110111: c <= 9'b1000110;
				8'b1011101: c <= 9'b1111;
				8'b1011011: c <= 9'b101001011;
				8'b111001: c <= 9'b100011000;
				8'b1001010: c <= 9'b1110010;
				8'b110011: c <= 9'b1111001;
				8'b1101100: c <= 9'b10111;
				8'b1110111: c <= 9'b101100101;
				8'b101011: c <= 9'b110111000;
				8'b1101011: c <= 9'b101110101;
				8'b111100: c <= 9'b10010110;
				8'b1000111: c <= 9'b110000;
				8'b1011111: c <= 9'b110111100;
				8'b1110100: c <= 9'b10100110;
				8'b101101: c <= 9'b111010100;
				8'b1010011: c <= 9'b11110100;
				8'b1100001: c <= 9'b110000001;
				8'b110101: c <= 9'b10010001;
				8'b1000100: c <= 9'b100;
				8'b1010001: c <= 9'b1111001;
				8'b1010100: c <= 9'b100111111;
				8'b1100110: c <= 9'b110001101;
				8'b101010: c <= 9'b1010110;
				8'b1011110: c <= 9'b110000010;
				8'b1100111: c <= 9'b11111100;
				8'b1011010: c <= 9'b101110111;
				8'b1000010: c <= 9'b101011010;
				8'b111101: c <= 9'b110111001;
				8'b110000: c <= 9'b110111;
				8'b111110: c <= 9'b1110;
				8'b1100010: c <= 9'b10111;
				8'b1110000: c <= 9'b11100010;
				8'b1101001: c <= 9'b1111001;
				8'b1110011: c <= 9'b10111001;
				8'b1001100: c <= 9'b101100000;
				8'b100001: c <= 9'b100011;
				8'b1000110: c <= 9'b110000010;
				8'b1110010: c <= 9'b111000101;
				8'b1010000: c <= 9'b100001;
				8'b1111010: c <= 9'b110010010;
				8'b1010101: c <= 9'b101011011;
				8'b111011: c <= 9'b101101100;
				8'b1001101: c <= 9'b110101100;
				8'b111111: c <= 9'b111000101;
				8'b1101110: c <= 9'b11011000;
				8'b1111011: c <= 9'b110111110;
				8'b1001011: c <= 9'b100110011;
				8'b1101111: c <= 9'b11000111;
				8'b1101000: c <= 9'b10101001;
				8'b101100: c <= 9'b1000000;
				8'b100100: c <= 9'b101010000;
				8'b1111000: c <= 9'b1010110;
				8'b1000101: c <= 9'b11011110;
				8'b1011001: c <= 9'b111101101;
				8'b110100: c <= 9'b101001;
				8'b1111001: c <= 9'b1001101;
				8'b1110001: c <= 9'b100100;
				8'b1001111: c <= 9'b11110;
				8'b1100101: c <= 9'b10001001;
				8'b1111110: c <= 9'b10111001;
				8'b1111100: c <= 9'b111010001;
				8'b1010110: c <= 9'b111111010;
				8'b110010: c <= 9'b111100010;
				8'b1101101: c <= 9'b111011111;
				8'b100011: c <= 9'b111011001;
				8'b1110101: c <= 9'b1010001;
				8'b1111101: c <= 9'b1111101;
				8'b101001: c <= 9'b1000101;
				8'b1010010: c <= 9'b10010011;
				8'b1011000: c <= 9'b10110010;
				8'b101110: c <= 9'b10001001;
				8'b1000001: c <= 9'b11010001;
				default: c <= 9'b0;
			endcase
			9'b111111111 : case(di)
				8'b1000011: c <= 9'b10101110;
				8'b101000: c <= 9'b10101100;
				8'b111010: c <= 9'b100011100;
				8'b110110: c <= 9'b111000101;
				8'b1100100: c <= 9'b101101001;
				8'b1000000: c <= 9'b11100;
				8'b1110110: c <= 9'b101100000;
				8'b100101: c <= 9'b100101;
				8'b101111: c <= 9'b101010;
				8'b100110: c <= 9'b10110110;
				8'b1100011: c <= 9'b110101110;
				8'b1001000: c <= 9'b11100111;
				8'b111000: c <= 9'b101000001;
				8'b110001: c <= 9'b1110;
				8'b1010111: c <= 9'b11010010;
				8'b1001110: c <= 9'b11000111;
				8'b1101010: c <= 9'b110011111;
				8'b1001001: c <= 9'b110011001;
				8'b1100000: c <= 9'b10111010;
				8'b110111: c <= 9'b10;
				8'b1011101: c <= 9'b110001;
				8'b1011011: c <= 9'b110000010;
				8'b111001: c <= 9'b100001111;
				8'b1001010: c <= 9'b10101011;
				8'b110011: c <= 9'b100010001;
				8'b1101100: c <= 9'b110101111;
				8'b1110111: c <= 9'b100100101;
				8'b101011: c <= 9'b111010100;
				8'b1101011: c <= 9'b100111100;
				8'b111100: c <= 9'b11101011;
				8'b1000111: c <= 9'b111100010;
				8'b1011111: c <= 9'b1100011;
				8'b1110100: c <= 9'b100010;
				8'b101101: c <= 9'b110110011;
				8'b1010011: c <= 9'b11100010;
				8'b1100001: c <= 9'b11001000;
				8'b110101: c <= 9'b100010100;
				8'b1000100: c <= 9'b111100111;
				8'b1010001: c <= 9'b110111000;
				8'b1010100: c <= 9'b1111;
				8'b1100110: c <= 9'b100001110;
				8'b101010: c <= 9'b101110110;
				8'b1011110: c <= 9'b10000001;
				8'b1100111: c <= 9'b100001111;
				8'b1011010: c <= 9'b111010100;
				8'b1000010: c <= 9'b11000100;
				8'b111101: c <= 9'b1110001;
				8'b110000: c <= 9'b110001;
				8'b111110: c <= 9'b100101010;
				8'b1100010: c <= 9'b100111000;
				8'b1110000: c <= 9'b101010110;
				8'b1101001: c <= 9'b10100010;
				8'b1110011: c <= 9'b10011011;
				8'b1001100: c <= 9'b111011100;
				8'b100001: c <= 9'b11111;
				8'b1000110: c <= 9'b110110000;
				8'b1110010: c <= 9'b1111010;
				8'b1010000: c <= 9'b101001010;
				8'b1111010: c <= 9'b1101101;
				8'b1010101: c <= 9'b111101000;
				8'b111011: c <= 9'b10110011;
				8'b1001101: c <= 9'b10000111;
				8'b111111: c <= 9'b11111;
				8'b1101110: c <= 9'b11101011;
				8'b1111011: c <= 9'b100111111;
				8'b1001011: c <= 9'b100000110;
				8'b1101111: c <= 9'b1100101;
				8'b1101000: c <= 9'b101001100;
				8'b101100: c <= 9'b110110010;
				8'b100100: c <= 9'b11000010;
				8'b1111000: c <= 9'b110110000;
				8'b1000101: c <= 9'b1110111;
				8'b1011001: c <= 9'b110100010;
				8'b110100: c <= 9'b101101010;
				8'b1111001: c <= 9'b111100110;
				8'b1110001: c <= 9'b11000000;
				8'b1001111: c <= 9'b100010111;
				8'b1100101: c <= 9'b10001100;
				8'b1111110: c <= 9'b10110100;
				8'b1111100: c <= 9'b111100101;
				8'b1010110: c <= 9'b1101101;
				8'b110010: c <= 9'b101011;
				8'b1101101: c <= 9'b101010110;
				8'b100011: c <= 9'b100011101;
				8'b1110101: c <= 9'b1001001;
				8'b1111101: c <= 9'b1001110;
				8'b101001: c <= 9'b111101110;
				8'b1010010: c <= 9'b10000011;
				8'b1011000: c <= 9'b1001010;
				8'b101110: c <= 9'b111011101;
				8'b1000001: c <= 9'b111100;
				default: c <= 9'b0;
			endcase
			9'b100011011 : case(di)
				8'b1000011: c <= 9'b101100011;
				8'b101000: c <= 9'b101011;
				8'b111010: c <= 9'b1110111;
				8'b110110: c <= 9'b101110100;
				8'b1100100: c <= 9'b100000111;
				8'b1000000: c <= 9'b10010101;
				8'b1110110: c <= 9'b101111010;
				8'b100101: c <= 9'b110001111;
				8'b101111: c <= 9'b100100001;
				8'b100110: c <= 9'b100110110;
				8'b1100011: c <= 9'b1110111;
				8'b1001000: c <= 9'b11110010;
				8'b111000: c <= 9'b11010101;
				8'b110001: c <= 9'b100011100;
				8'b1010111: c <= 9'b1111100;
				8'b1001110: c <= 9'b11100110;
				8'b1101010: c <= 9'b111001;
				8'b1001001: c <= 9'b10101110;
				8'b1100000: c <= 9'b11101011;
				8'b110111: c <= 9'b10011010;
				8'b1011101: c <= 9'b101010101;
				8'b1011011: c <= 9'b101000110;
				8'b111001: c <= 9'b10000;
				8'b1001010: c <= 9'b10100101;
				8'b110011: c <= 9'b101111001;
				8'b1101100: c <= 9'b111111;
				8'b1110111: c <= 9'b100000011;
				8'b101011: c <= 9'b11011110;
				8'b1101011: c <= 9'b10011010;
				8'b111100: c <= 9'b11001001;
				8'b1000111: c <= 9'b111011100;
				8'b1011111: c <= 9'b11011100;
				8'b1110100: c <= 9'b11000000;
				8'b101101: c <= 9'b11110111;
				8'b1010011: c <= 9'b110101101;
				8'b1100001: c <= 9'b101000;
				8'b110101: c <= 9'b10111;
				8'b1000100: c <= 9'b100110000;
				8'b1010001: c <= 9'b110001001;
				8'b1010100: c <= 9'b11110110;
				8'b1100110: c <= 9'b101101101;
				8'b101010: c <= 9'b110101100;
				8'b1011110: c <= 9'b1111111;
				8'b1100111: c <= 9'b1000011;
				8'b1011010: c <= 9'b110010100;
				8'b1000010: c <= 9'b100110110;
				8'b111101: c <= 9'b111010000;
				8'b110000: c <= 9'b101101100;
				8'b111110: c <= 9'b110100111;
				8'b1100010: c <= 9'b110110;
				8'b1110000: c <= 9'b111001110;
				8'b1101001: c <= 9'b101111010;
				8'b1110011: c <= 9'b10110100;
				8'b1001100: c <= 9'b110000101;
				8'b100001: c <= 9'b110011011;
				8'b1000110: c <= 9'b1000;
				8'b1110010: c <= 9'b10100110;
				8'b1010000: c <= 9'b110101010;
				8'b1111010: c <= 9'b1100011;
				8'b1010101: c <= 9'b111110001;
				8'b111011: c <= 9'b1010011;
				8'b1001101: c <= 9'b110100101;
				8'b111111: c <= 9'b11011000;
				8'b1101110: c <= 9'b1111001;
				8'b1111011: c <= 9'b1000101;
				8'b1001011: c <= 9'b110101011;
				8'b1101111: c <= 9'b10101110;
				8'b1101000: c <= 9'b100100001;
				8'b101100: c <= 9'b10011101;
				8'b100100: c <= 9'b110001010;
				8'b1111000: c <= 9'b111000000;
				8'b1000101: c <= 9'b11011101;
				8'b1011001: c <= 9'b101111110;
				8'b110100: c <= 9'b11011011;
				8'b1111001: c <= 9'b1101010;
				8'b1110001: c <= 9'b10111111;
				8'b1001111: c <= 9'b10111110;
				8'b1100101: c <= 9'b1100;
				8'b1111110: c <= 9'b10101111;
				8'b1111100: c <= 9'b11111000;
				8'b1010110: c <= 9'b111100011;
				8'b110010: c <= 9'b1110000;
				8'b1101101: c <= 9'b110011;
				8'b100011: c <= 9'b110010101;
				8'b1110101: c <= 9'b100010110;
				8'b1111101: c <= 9'b101011101;
				8'b101001: c <= 9'b11111001;
				8'b1010010: c <= 9'b1001000;
				8'b1011000: c <= 9'b101001000;
				8'b101110: c <= 9'b11000;
				8'b1000001: c <= 9'b10110001;
				default: c <= 9'b0;
			endcase
			9'b110000000 : case(di)
				8'b1000011: c <= 9'b100100110;
				8'b101000: c <= 9'b111110110;
				8'b111010: c <= 9'b1110111;
				8'b110110: c <= 9'b11110001;
				8'b1100100: c <= 9'b110001;
				8'b1000000: c <= 9'b10000101;
				8'b1110110: c <= 9'b11101111;
				8'b100101: c <= 9'b110011010;
				8'b101111: c <= 9'b1100111;
				8'b100110: c <= 9'b100010011;
				8'b1100011: c <= 9'b1001001;
				8'b1001000: c <= 9'b1111011;
				8'b111000: c <= 9'b11011001;
				8'b110001: c <= 9'b1011100;
				8'b1010111: c <= 9'b100010001;
				8'b1001110: c <= 9'b110100111;
				8'b1101010: c <= 9'b11001010;
				8'b1001001: c <= 9'b10101000;
				8'b1100000: c <= 9'b100011100;
				8'b110111: c <= 9'b10101010;
				8'b1011101: c <= 9'b101010000;
				8'b1011011: c <= 9'b11110101;
				8'b111001: c <= 9'b101101110;
				8'b1001010: c <= 9'b10000110;
				8'b110011: c <= 9'b10100111;
				8'b1101100: c <= 9'b100011000;
				8'b1110111: c <= 9'b11010101;
				8'b101011: c <= 9'b111010100;
				8'b1101011: c <= 9'b110100110;
				8'b111100: c <= 9'b11;
				8'b1000111: c <= 9'b100111;
				8'b1011111: c <= 9'b10000111;
				8'b1110100: c <= 9'b11100011;
				8'b101101: c <= 9'b110001011;
				8'b1010011: c <= 9'b11001111;
				8'b1100001: c <= 9'b101011011;
				8'b110101: c <= 9'b110001010;
				8'b1000100: c <= 9'b110110100;
				8'b1010001: c <= 9'b111001010;
				8'b1010100: c <= 9'b1111000;
				8'b1100110: c <= 9'b10110010;
				8'b101010: c <= 9'b110010011;
				8'b1011110: c <= 9'b10010011;
				8'b1100111: c <= 9'b100001001;
				8'b1011010: c <= 9'b111101;
				8'b1000010: c <= 9'b100011100;
				8'b111101: c <= 9'b11110;
				8'b110000: c <= 9'b1101110;
				8'b111110: c <= 9'b1001000;
				8'b1100010: c <= 9'b100010011;
				8'b1110000: c <= 9'b101101011;
				8'b1101001: c <= 9'b1011100;
				8'b1110011: c <= 9'b101011101;
				8'b1001100: c <= 9'b101001011;
				8'b100001: c <= 9'b10111111;
				8'b1000110: c <= 9'b10100010;
				8'b1110010: c <= 9'b101010000;
				8'b1010000: c <= 9'b111111011;
				8'b1111010: c <= 9'b100010;
				8'b1010101: c <= 9'b100110010;
				8'b111011: c <= 9'b1001111;
				8'b1001101: c <= 9'b10000111;
				8'b111111: c <= 9'b1000101;
				8'b1101110: c <= 9'b10100111;
				8'b1111011: c <= 9'b100000100;
				8'b1001011: c <= 9'b11101100;
				8'b1101111: c <= 9'b110000111;
				8'b1101000: c <= 9'b10111111;
				8'b101100: c <= 9'b111010000;
				8'b100100: c <= 9'b101110100;
				8'b1111000: c <= 9'b101011011;
				8'b1000101: c <= 9'b101100100;
				8'b1011001: c <= 9'b101001000;
				8'b110100: c <= 9'b10010100;
				8'b1111001: c <= 9'b1001101;
				8'b1110001: c <= 9'b101110111;
				8'b1001111: c <= 9'b10111001;
				8'b1100101: c <= 9'b100011001;
				8'b1111110: c <= 9'b100;
				8'b1111100: c <= 9'b111111010;
				8'b1010110: c <= 9'b101010111;
				8'b110010: c <= 9'b111111001;
				8'b1101101: c <= 9'b100101001;
				8'b100011: c <= 9'b1110001;
				8'b1110101: c <= 9'b110000111;
				8'b1111101: c <= 9'b110101101;
				8'b101001: c <= 9'b110000010;
				8'b1010010: c <= 9'b110011101;
				8'b1011000: c <= 9'b1000101;
				8'b101110: c <= 9'b111010000;
				8'b1000001: c <= 9'b1001010;
				default: c <= 9'b0;
			endcase
			9'b11011101 : case(di)
				8'b1000011: c <= 9'b111011111;
				8'b101000: c <= 9'b101110001;
				8'b111010: c <= 9'b111101;
				8'b110110: c <= 9'b100100010;
				8'b1100100: c <= 9'b11100011;
				8'b1000000: c <= 9'b100000111;
				8'b1110110: c <= 9'b10001011;
				8'b100101: c <= 9'b100010010;
				8'b101111: c <= 9'b10011001;
				8'b100110: c <= 9'b110010;
				8'b1100011: c <= 9'b10011011;
				8'b1001000: c <= 9'b11000110;
				8'b111000: c <= 9'b100010000;
				8'b110001: c <= 9'b1101000;
				8'b1010111: c <= 9'b110110110;
				8'b1001110: c <= 9'b110101110;
				8'b1101010: c <= 9'b101011001;
				8'b1001001: c <= 9'b1001001;
				8'b1100000: c <= 9'b1111001;
				8'b110111: c <= 9'b110100111;
				8'b1011101: c <= 9'b1010010;
				8'b1011011: c <= 9'b100111001;
				8'b111001: c <= 9'b11001;
				8'b1001010: c <= 9'b10110100;
				8'b110011: c <= 9'b10110010;
				8'b1101100: c <= 9'b100110101;
				8'b1110111: c <= 9'b110100010;
				8'b101011: c <= 9'b111000100;
				8'b1101011: c <= 9'b10100010;
				8'b111100: c <= 9'b100101101;
				8'b1000111: c <= 9'b11110000;
				8'b1011111: c <= 9'b100100011;
				8'b1110100: c <= 9'b101110100;
				8'b101101: c <= 9'b11000000;
				8'b1010011: c <= 9'b11100110;
				8'b1100001: c <= 9'b1000011;
				8'b110101: c <= 9'b1101000;
				8'b1000100: c <= 9'b1001;
				8'b1010001: c <= 9'b101000011;
				8'b1010100: c <= 9'b110010101;
				8'b1100110: c <= 9'b101100010;
				8'b101010: c <= 9'b111100;
				8'b1011110: c <= 9'b110111110;
				8'b1100111: c <= 9'b101011001;
				8'b1011010: c <= 9'b111011111;
				8'b1000010: c <= 9'b101010101;
				8'b111101: c <= 9'b11111;
				8'b110000: c <= 9'b10001000;
				8'b111110: c <= 9'b111101010;
				8'b1100010: c <= 9'b10111010;
				8'b1110000: c <= 9'b110100;
				8'b1101001: c <= 9'b10000101;
				8'b1110011: c <= 9'b10010000;
				8'b1001100: c <= 9'b110101110;
				8'b100001: c <= 9'b110001111;
				8'b1000110: c <= 9'b1110010;
				8'b1110010: c <= 9'b111101110;
				8'b1010000: c <= 9'b1101110;
				8'b1111010: c <= 9'b101110;
				8'b1010101: c <= 9'b1100011;
				8'b111011: c <= 9'b11100;
				8'b1001101: c <= 9'b101100100;
				8'b111111: c <= 9'b11000111;
				8'b1101110: c <= 9'b110001111;
				8'b1111011: c <= 9'b101111010;
				8'b1001011: c <= 9'b110001000;
				8'b1101111: c <= 9'b10000110;
				8'b1101000: c <= 9'b111110110;
				8'b101100: c <= 9'b1;
				8'b100100: c <= 9'b101011000;
				8'b1111000: c <= 9'b11100110;
				8'b1000101: c <= 9'b11010101;
				8'b1011001: c <= 9'b10011100;
				8'b110100: c <= 9'b1011010;
				8'b1111001: c <= 9'b10011010;
				8'b1110001: c <= 9'b100101111;
				8'b1001111: c <= 9'b1000101;
				8'b1100101: c <= 9'b111001101;
				8'b1111110: c <= 9'b1001001;
				8'b1111100: c <= 9'b11001111;
				8'b1010110: c <= 9'b111100001;
				8'b110010: c <= 9'b101001100;
				8'b1101101: c <= 9'b110011011;
				8'b100011: c <= 9'b110001;
				8'b1110101: c <= 9'b10001111;
				8'b1111101: c <= 9'b11001001;
				8'b101001: c <= 9'b101000;
				8'b1010010: c <= 9'b100101011;
				8'b1011000: c <= 9'b101100000;
				8'b101110: c <= 9'b1000110;
				8'b1000001: c <= 9'b11000010;
				default: c <= 9'b0;
			endcase
			9'b11000110 : case(di)
				8'b1000011: c <= 9'b101101110;
				8'b101000: c <= 9'b100001011;
				8'b111010: c <= 9'b100100001;
				8'b110110: c <= 9'b111010001;
				8'b1100100: c <= 9'b10101110;
				8'b1000000: c <= 9'b100101100;
				8'b1110110: c <= 9'b11100100;
				8'b100101: c <= 9'b110011111;
				8'b101111: c <= 9'b1000101;
				8'b100110: c <= 9'b1001010;
				8'b1100011: c <= 9'b100110000;
				8'b1001000: c <= 9'b11101011;
				8'b111000: c <= 9'b10000000;
				8'b110001: c <= 9'b10001101;
				8'b1010111: c <= 9'b10100110;
				8'b1001110: c <= 9'b111001111;
				8'b1101010: c <= 9'b10110;
				8'b1001001: c <= 9'b11001;
				8'b1100000: c <= 9'b11010011;
				8'b110111: c <= 9'b101100111;
				8'b1011101: c <= 9'b11111;
				8'b1011011: c <= 9'b111001011;
				8'b111001: c <= 9'b101001000;
				8'b1001010: c <= 9'b110010110;
				8'b110011: c <= 9'b101111110;
				8'b1101100: c <= 9'b1101111;
				8'b1110111: c <= 9'b11100100;
				8'b101011: c <= 9'b11101;
				8'b1101011: c <= 9'b100110111;
				8'b111100: c <= 9'b110100010;
				8'b1000111: c <= 9'b111100010;
				8'b1011111: c <= 9'b1110010;
				8'b1110100: c <= 9'b111101010;
				8'b101101: c <= 9'b10100011;
				8'b1010011: c <= 9'b111;
				8'b1100001: c <= 9'b111100111;
				8'b110101: c <= 9'b11101100;
				8'b1000100: c <= 9'b11010100;
				8'b1010001: c <= 9'b10100000;
				8'b1010100: c <= 9'b111000110;
				8'b1100110: c <= 9'b111001011;
				8'b101010: c <= 9'b101101;
				8'b1011110: c <= 9'b100100011;
				8'b1100111: c <= 9'b111110110;
				8'b1011010: c <= 9'b110110100;
				8'b1000010: c <= 9'b110100011;
				8'b111101: c <= 9'b10000000;
				8'b110000: c <= 9'b11111001;
				8'b111110: c <= 9'b1011001;
				8'b1100010: c <= 9'b10001110;
				8'b1110000: c <= 9'b1111001;
				8'b1101001: c <= 9'b110010101;
				8'b1110011: c <= 9'b111110101;
				8'b1001100: c <= 9'b10001101;
				8'b100001: c <= 9'b100001001;
				8'b1000110: c <= 9'b1000011;
				8'b1110010: c <= 9'b10111111;
				8'b1010000: c <= 9'b100000100;
				8'b1111010: c <= 9'b110011001;
				8'b1010101: c <= 9'b100111101;
				8'b111011: c <= 9'b10001011;
				8'b1001101: c <= 9'b1111;
				8'b111111: c <= 9'b100110010;
				8'b1101110: c <= 9'b10000;
				8'b1111011: c <= 9'b1001000;
				8'b1001011: c <= 9'b100110010;
				8'b1101111: c <= 9'b100001111;
				8'b1101000: c <= 9'b10010;
				8'b101100: c <= 9'b111001110;
				8'b100100: c <= 9'b11100010;
				8'b1111000: c <= 9'b10110111;
				8'b1000101: c <= 9'b10011011;
				8'b1011001: c <= 9'b111111;
				8'b110100: c <= 9'b1000001;
				8'b1111001: c <= 9'b100101001;
				8'b1110001: c <= 9'b101010;
				8'b1001111: c <= 9'b10001010;
				8'b1100101: c <= 9'b110110010;
				8'b1111110: c <= 9'b11110101;
				8'b1111100: c <= 9'b1101;
				8'b1010110: c <= 9'b10000000;
				8'b110010: c <= 9'b101101100;
				8'b1101101: c <= 9'b1000000;
				8'b100011: c <= 9'b100101010;
				8'b1110101: c <= 9'b101001000;
				8'b1111101: c <= 9'b101001010;
				8'b101001: c <= 9'b100010100;
				8'b1010010: c <= 9'b10111001;
				8'b1011000: c <= 9'b100001;
				8'b101110: c <= 9'b101001110;
				8'b1000001: c <= 9'b10110011;
				default: c <= 9'b0;
			endcase
			9'b100010011 : case(di)
				8'b1000011: c <= 9'b10110110;
				8'b101000: c <= 9'b11010101;
				8'b111010: c <= 9'b10110110;
				8'b110110: c <= 9'b100001001;
				8'b1100100: c <= 9'b111010100;
				8'b1000000: c <= 9'b100111011;
				8'b1110110: c <= 9'b100001;
				8'b100101: c <= 9'b10000101;
				8'b101111: c <= 9'b110101001;
				8'b100110: c <= 9'b1100100;
				8'b1100011: c <= 9'b10100011;
				8'b1001000: c <= 9'b110011;
				8'b111000: c <= 9'b10101110;
				8'b110001: c <= 9'b101100000;
				8'b1010111: c <= 9'b10000101;
				8'b1001110: c <= 9'b100001101;
				8'b1101010: c <= 9'b101010011;
				8'b1001001: c <= 9'b110111001;
				8'b1100000: c <= 9'b100101100;
				8'b110111: c <= 9'b110101101;
				8'b1011101: c <= 9'b10000010;
				8'b1011011: c <= 9'b111100101;
				8'b111001: c <= 9'b100110;
				8'b1001010: c <= 9'b1110101;
				8'b110011: c <= 9'b111001011;
				8'b1101100: c <= 9'b100011111;
				8'b1110111: c <= 9'b101010001;
				8'b101011: c <= 9'b1010001;
				8'b1101011: c <= 9'b10100;
				8'b111100: c <= 9'b1011010;
				8'b1000111: c <= 9'b1101110;
				8'b1011111: c <= 9'b100001010;
				8'b1110100: c <= 9'b101110111;
				8'b101101: c <= 9'b1100000;
				8'b1010011: c <= 9'b101;
				8'b1100001: c <= 9'b110000000;
				8'b110101: c <= 9'b110000001;
				8'b1000100: c <= 9'b111101000;
				8'b1010001: c <= 9'b10011;
				8'b1010100: c <= 9'b110011111;
				8'b1100110: c <= 9'b101000111;
				8'b101010: c <= 9'b10101010;
				8'b1011110: c <= 9'b101110111;
				8'b1100111: c <= 9'b111100011;
				8'b1011010: c <= 9'b10011011;
				8'b1000010: c <= 9'b110100011;
				8'b111101: c <= 9'b1011;
				8'b110000: c <= 9'b1010011;
				8'b111110: c <= 9'b110010101;
				8'b1100010: c <= 9'b11001;
				8'b1110000: c <= 9'b1100100;
				8'b1101001: c <= 9'b100010001;
				8'b1110011: c <= 9'b101100101;
				8'b1001100: c <= 9'b11111101;
				8'b100001: c <= 9'b101011001;
				8'b1000110: c <= 9'b1011;
				8'b1110010: c <= 9'b111111110;
				8'b1010000: c <= 9'b111010000;
				8'b1111010: c <= 9'b100101010;
				8'b1010101: c <= 9'b11001001;
				8'b111011: c <= 9'b110001011;
				8'b1001101: c <= 9'b100010101;
				8'b111111: c <= 9'b100111110;
				8'b1101110: c <= 9'b111011100;
				8'b1111011: c <= 9'b1001;
				8'b1001011: c <= 9'b1110100;
				8'b1101111: c <= 9'b111001;
				8'b1101000: c <= 9'b111101;
				8'b101100: c <= 9'b101101000;
				8'b100100: c <= 9'b110010100;
				8'b1111000: c <= 9'b11111;
				8'b1000101: c <= 9'b11001110;
				8'b1011001: c <= 9'b11010101;
				8'b110100: c <= 9'b1110111;
				8'b1111001: c <= 9'b101101;
				8'b1110001: c <= 9'b101010001;
				8'b1001111: c <= 9'b111101110;
				8'b1100101: c <= 9'b1110011;
				8'b1111110: c <= 9'b101010101;
				8'b1111100: c <= 9'b101110010;
				8'b1010110: c <= 9'b10101001;
				8'b110010: c <= 9'b101111000;
				8'b1101101: c <= 9'b10011;
				8'b100011: c <= 9'b11000000;
				8'b1110101: c <= 9'b111011;
				8'b1111101: c <= 9'b1010111;
				8'b101001: c <= 9'b10001010;
				8'b1010010: c <= 9'b11110;
				8'b1011000: c <= 9'b101101;
				8'b101110: c <= 9'b100100011;
				8'b1000001: c <= 9'b100110000;
				default: c <= 9'b0;
			endcase
			9'b111101010 : case(di)
				8'b1000011: c <= 9'b11010000;
				8'b101000: c <= 9'b101000;
				8'b111010: c <= 9'b110001001;
				8'b110110: c <= 9'b111011011;
				8'b1100100: c <= 9'b101000001;
				8'b1000000: c <= 9'b1101110;
				8'b1110110: c <= 9'b100011011;
				8'b100101: c <= 9'b110101011;
				8'b101111: c <= 9'b10110001;
				8'b100110: c <= 9'b101101;
				8'b1100011: c <= 9'b1100001;
				8'b1001000: c <= 9'b101111110;
				8'b111000: c <= 9'b10111;
				8'b110001: c <= 9'b101100101;
				8'b1010111: c <= 9'b11010100;
				8'b1001110: c <= 9'b100111;
				8'b1101010: c <= 9'b100001101;
				8'b1001001: c <= 9'b111101;
				8'b1100000: c <= 9'b101110100;
				8'b110111: c <= 9'b100001001;
				8'b1011101: c <= 9'b111100100;
				8'b1011011: c <= 9'b111100100;
				8'b111001: c <= 9'b11100000;
				8'b1001010: c <= 9'b100100101;
				8'b110011: c <= 9'b101010100;
				8'b1101100: c <= 9'b100101100;
				8'b1110111: c <= 9'b110000000;
				8'b101011: c <= 9'b110001001;
				8'b1101011: c <= 9'b111001101;
				8'b111100: c <= 9'b100011001;
				8'b1000111: c <= 9'b100010000;
				8'b1011111: c <= 9'b100000101;
				8'b1110100: c <= 9'b100101000;
				8'b101101: c <= 9'b110100101;
				8'b1010011: c <= 9'b1101000;
				8'b1100001: c <= 9'b111001101;
				8'b110101: c <= 9'b110100101;
				8'b1000100: c <= 9'b10101;
				8'b1010001: c <= 9'b110110110;
				8'b1010100: c <= 9'b110010001;
				8'b1100110: c <= 9'b100001010;
				8'b101010: c <= 9'b10011101;
				8'b1011110: c <= 9'b10100;
				8'b1100111: c <= 9'b11110100;
				8'b1011010: c <= 9'b10101000;
				8'b1000010: c <= 9'b10100011;
				8'b111101: c <= 9'b11101101;
				8'b110000: c <= 9'b110100101;
				8'b111110: c <= 9'b100000011;
				8'b1100010: c <= 9'b11000000;
				8'b1110000: c <= 9'b111011111;
				8'b1101001: c <= 9'b100010011;
				8'b1110011: c <= 9'b111101;
				8'b1001100: c <= 9'b1110111;
				8'b100001: c <= 9'b111111101;
				8'b1000110: c <= 9'b11011110;
				8'b1110010: c <= 9'b100110000;
				8'b1010000: c <= 9'b101000010;
				8'b1111010: c <= 9'b1010000;
				8'b1010101: c <= 9'b101001100;
				8'b111011: c <= 9'b111000100;
				8'b1001101: c <= 9'b100110111;
				8'b111111: c <= 9'b1011011;
				8'b1101110: c <= 9'b10001010;
				8'b1111011: c <= 9'b101011001;
				8'b1001011: c <= 9'b11101100;
				8'b1101111: c <= 9'b110110010;
				8'b1101000: c <= 9'b110100111;
				8'b101100: c <= 9'b10010100;
				8'b100100: c <= 9'b10101;
				8'b1111000: c <= 9'b1110101;
				8'b1000101: c <= 9'b110110011;
				8'b1011001: c <= 9'b111001101;
				8'b110100: c <= 9'b11010111;
				8'b1111001: c <= 9'b101110101;
				8'b1110001: c <= 9'b101101;
				8'b1001111: c <= 9'b10101101;
				8'b1100101: c <= 9'b111100;
				8'b1111110: c <= 9'b11110101;
				8'b1111100: c <= 9'b110000000;
				8'b1010110: c <= 9'b100011;
				8'b110010: c <= 9'b1010111;
				8'b1101101: c <= 9'b111110110;
				8'b100011: c <= 9'b1011100;
				8'b1110101: c <= 9'b11;
				8'b1111101: c <= 9'b100100;
				8'b101001: c <= 9'b111100010;
				8'b1010010: c <= 9'b110000010;
				8'b1011000: c <= 9'b110010110;
				8'b101110: c <= 9'b100001111;
				8'b1000001: c <= 9'b1100000;
				default: c <= 9'b0;
			endcase
			9'b100011111 : case(di)
				8'b1000011: c <= 9'b100111010;
				8'b101000: c <= 9'b1000100;
				8'b111010: c <= 9'b10100010;
				8'b110110: c <= 9'b10011100;
				8'b1100100: c <= 9'b101101101;
				8'b1000000: c <= 9'b101110100;
				8'b1110110: c <= 9'b100101010;
				8'b100101: c <= 9'b11101111;
				8'b101111: c <= 9'b1000000;
				8'b100110: c <= 9'b1000011;
				8'b1100011: c <= 9'b1011000;
				8'b1001000: c <= 9'b111111111;
				8'b111000: c <= 9'b111111;
				8'b110001: c <= 9'b11000;
				8'b1010111: c <= 9'b10010;
				8'b1001110: c <= 9'b11111011;
				8'b1101010: c <= 9'b101100101;
				8'b1001001: c <= 9'b11000100;
				8'b1100000: c <= 9'b10111;
				8'b110111: c <= 9'b10100000;
				8'b1011101: c <= 9'b10001000;
				8'b1011011: c <= 9'b111110000;
				8'b111001: c <= 9'b101111111;
				8'b1001010: c <= 9'b10000101;
				8'b110011: c <= 9'b10011111;
				8'b1101100: c <= 9'b110011010;
				8'b1110111: c <= 9'b101100111;
				8'b101011: c <= 9'b110101100;
				8'b1101011: c <= 9'b11010010;
				8'b111100: c <= 9'b1111011;
				8'b1000111: c <= 9'b10011000;
				8'b1011111: c <= 9'b110;
				8'b1110100: c <= 9'b10000110;
				8'b101101: c <= 9'b100101110;
				8'b1010011: c <= 9'b111101101;
				8'b1100001: c <= 9'b1000000;
				8'b110101: c <= 9'b11011100;
				8'b1000100: c <= 9'b101010111;
				8'b1010001: c <= 9'b100111111;
				8'b1010100: c <= 9'b1001011;
				8'b1100110: c <= 9'b1001;
				8'b101010: c <= 9'b100011010;
				8'b1011110: c <= 9'b11110011;
				8'b1100111: c <= 9'b100110011;
				8'b1011010: c <= 9'b1001111;
				8'b1000010: c <= 9'b110011110;
				8'b111101: c <= 9'b1111;
				8'b110000: c <= 9'b110000;
				8'b111110: c <= 9'b100111110;
				8'b1100010: c <= 9'b1000101;
				8'b1110000: c <= 9'b110011110;
				8'b1101001: c <= 9'b111101;
				8'b1110011: c <= 9'b11001101;
				8'b1001100: c <= 9'b10111001;
				8'b100001: c <= 9'b111100110;
				8'b1000110: c <= 9'b111000100;
				8'b1110010: c <= 9'b111011010;
				8'b1010000: c <= 9'b101101001;
				8'b1111010: c <= 9'b111001000;
				8'b1010101: c <= 9'b110110101;
				8'b111011: c <= 9'b1011110;
				8'b1001101: c <= 9'b100101011;
				8'b111111: c <= 9'b1001011;
				8'b1101110: c <= 9'b10110001;
				8'b1111011: c <= 9'b1110101;
				8'b1001011: c <= 9'b11011010;
				8'b1101111: c <= 9'b11010111;
				8'b1101000: c <= 9'b101010011;
				8'b101100: c <= 9'b1001000;
				8'b100100: c <= 9'b10101101;
				8'b1111000: c <= 9'b110001100;
				8'b1000101: c <= 9'b111110001;
				8'b1011001: c <= 9'b100001;
				8'b110100: c <= 9'b110011100;
				8'b1111001: c <= 9'b10011000;
				8'b1110001: c <= 9'b11100010;
				8'b1001111: c <= 9'b110011110;
				8'b1100101: c <= 9'b11100110;
				8'b1111110: c <= 9'b101001100;
				8'b1111100: c <= 9'b111001010;
				8'b1010110: c <= 9'b110110111;
				8'b110010: c <= 9'b101100100;
				8'b1101101: c <= 9'b1101010;
				8'b100011: c <= 9'b110011010;
				8'b1110101: c <= 9'b1101010;
				8'b1111101: c <= 9'b111100100;
				8'b101001: c <= 9'b11110010;
				8'b1010010: c <= 9'b101000100;
				8'b1011000: c <= 9'b10001101;
				8'b101110: c <= 9'b101001010;
				8'b1000001: c <= 9'b100111001;
				default: c <= 9'b0;
			endcase
			9'b101100101 : case(di)
				8'b1000011: c <= 9'b101000011;
				8'b101000: c <= 9'b11100000;
				8'b111010: c <= 9'b100000011;
				8'b110110: c <= 9'b10101010;
				8'b1100100: c <= 9'b10001011;
				8'b1000000: c <= 9'b111000;
				8'b1110110: c <= 9'b10000101;
				8'b100101: c <= 9'b111001011;
				8'b101111: c <= 9'b10011;
				8'b100110: c <= 9'b110001001;
				8'b1100011: c <= 9'b101001001;
				8'b1001000: c <= 9'b101100111;
				8'b111000: c <= 9'b1101001;
				8'b110001: c <= 9'b11111100;
				8'b1010111: c <= 9'b110111;
				8'b1001110: c <= 9'b1000;
				8'b1101010: c <= 9'b110010010;
				8'b1001001: c <= 9'b100000000;
				8'b1100000: c <= 9'b1110111;
				8'b110111: c <= 9'b10000000;
				8'b1011101: c <= 9'b1010010;
				8'b1011011: c <= 9'b100100110;
				8'b111001: c <= 9'b101101110;
				8'b1001010: c <= 9'b110010101;
				8'b110011: c <= 9'b101111010;
				8'b1101100: c <= 9'b101100111;
				8'b1110111: c <= 9'b1011011;
				8'b101011: c <= 9'b10000000;
				8'b1101011: c <= 9'b101000111;
				8'b111100: c <= 9'b101111000;
				8'b1000111: c <= 9'b100110010;
				8'b1011111: c <= 9'b1100011;
				8'b1110100: c <= 9'b11001000;
				8'b101101: c <= 9'b100111101;
				8'b1010011: c <= 9'b110001001;
				8'b1100001: c <= 9'b10010101;
				8'b110101: c <= 9'b101000010;
				8'b1000100: c <= 9'b1000;
				8'b1010001: c <= 9'b100010100;
				8'b1010100: c <= 9'b11010101;
				8'b1100110: c <= 9'b111011110;
				8'b101010: c <= 9'b11100;
				8'b1011110: c <= 9'b101010011;
				8'b1100111: c <= 9'b10010011;
				8'b1011010: c <= 9'b10110111;
				8'b1000010: c <= 9'b101001000;
				8'b111101: c <= 9'b10000111;
				8'b110000: c <= 9'b100100010;
				8'b111110: c <= 9'b1000101;
				8'b1100010: c <= 9'b10100;
				8'b1110000: c <= 9'b10100000;
				8'b1101001: c <= 9'b1001100;
				8'b1110011: c <= 9'b110111011;
				8'b1001100: c <= 9'b1000110;
				8'b100001: c <= 9'b111000011;
				8'b1000110: c <= 9'b11111100;
				8'b1110010: c <= 9'b11000010;
				8'b1010000: c <= 9'b110101110;
				8'b1111010: c <= 9'b101001010;
				8'b1010101: c <= 9'b101001011;
				8'b111011: c <= 9'b110000001;
				8'b1001101: c <= 9'b11111;
				8'b111111: c <= 9'b110101011;
				8'b1101110: c <= 9'b10001011;
				8'b1111011: c <= 9'b111000;
				8'b1001011: c <= 9'b1000001;
				8'b1101111: c <= 9'b100100010;
				8'b1101000: c <= 9'b1000101;
				8'b101100: c <= 9'b101010;
				8'b100100: c <= 9'b101100011;
				8'b1111000: c <= 9'b101000011;
				8'b1000101: c <= 9'b100110010;
				8'b1011001: c <= 9'b1010101;
				8'b110100: c <= 9'b101001100;
				8'b1111001: c <= 9'b110100101;
				8'b1110001: c <= 9'b100000110;
				8'b1001111: c <= 9'b10100110;
				8'b1100101: c <= 9'b111000111;
				8'b1111110: c <= 9'b101001100;
				8'b1111100: c <= 9'b110101100;
				8'b1010110: c <= 9'b11010;
				8'b110010: c <= 9'b101000;
				8'b1101101: c <= 9'b100010000;
				8'b100011: c <= 9'b111001001;
				8'b1110101: c <= 9'b1100100;
				8'b1111101: c <= 9'b11100010;
				8'b101001: c <= 9'b101000011;
				8'b1010010: c <= 9'b1111010;
				8'b1011000: c <= 9'b110001011;
				8'b101110: c <= 9'b1100001;
				8'b1000001: c <= 9'b11110001;
				default: c <= 9'b0;
			endcase
			9'b11010111 : case(di)
				8'b1000011: c <= 9'b101100110;
				8'b101000: c <= 9'b1111110;
				8'b111010: c <= 9'b10011;
				8'b110110: c <= 9'b1111011;
				8'b1100100: c <= 9'b100101110;
				8'b1000000: c <= 9'b101101110;
				8'b1110110: c <= 9'b1001011;
				8'b100101: c <= 9'b11011010;
				8'b101111: c <= 9'b100111001;
				8'b100110: c <= 9'b101001100;
				8'b1100011: c <= 9'b11001010;
				8'b1001000: c <= 9'b110010001;
				8'b111000: c <= 9'b1111000;
				8'b110001: c <= 9'b111011011;
				8'b1010111: c <= 9'b100000001;
				8'b1001110: c <= 9'b111001011;
				8'b1101010: c <= 9'b100011000;
				8'b1001001: c <= 9'b110010101;
				8'b1100000: c <= 9'b10011101;
				8'b110111: c <= 9'b11010;
				8'b1011101: c <= 9'b1101100;
				8'b1011011: c <= 9'b101110110;
				8'b111001: c <= 9'b10111100;
				8'b1001010: c <= 9'b10011100;
				8'b110011: c <= 9'b101101011;
				8'b1101100: c <= 9'b101001110;
				8'b1110111: c <= 9'b1100000;
				8'b101011: c <= 9'b111001001;
				8'b1101011: c <= 9'b101100000;
				8'b111100: c <= 9'b100010111;
				8'b1000111: c <= 9'b110110101;
				8'b1011111: c <= 9'b11000010;
				8'b1110100: c <= 9'b111000110;
				8'b101101: c <= 9'b110000010;
				8'b1010011: c <= 9'b101000011;
				8'b1100001: c <= 9'b100010001;
				8'b110101: c <= 9'b11100;
				8'b1000100: c <= 9'b1010011;
				8'b1010001: c <= 9'b101110001;
				8'b1010100: c <= 9'b1110;
				8'b1100110: c <= 9'b110010101;
				8'b101010: c <= 9'b11010001;
				8'b1011110: c <= 9'b10011010;
				8'b1100111: c <= 9'b11100010;
				8'b1011010: c <= 9'b1100010;
				8'b1000010: c <= 9'b1000;
				8'b111101: c <= 9'b111000;
				8'b110000: c <= 9'b100000010;
				8'b111110: c <= 9'b111111010;
				8'b1100010: c <= 9'b10100;
				8'b1110000: c <= 9'b110111001;
				8'b1101001: c <= 9'b100010001;
				8'b1110011: c <= 9'b101101111;
				8'b1001100: c <= 9'b110001000;
				8'b100001: c <= 9'b100011011;
				8'b1000110: c <= 9'b101100101;
				8'b1110010: c <= 9'b1111011;
				8'b1010000: c <= 9'b111001101;
				8'b1111010: c <= 9'b10100111;
				8'b1010101: c <= 9'b101100111;
				8'b111011: c <= 9'b111001110;
				8'b1001101: c <= 9'b111101101;
				8'b111111: c <= 9'b111101;
				8'b1101110: c <= 9'b111111001;
				8'b1111011: c <= 9'b110101100;
				8'b1001011: c <= 9'b110110101;
				8'b1101111: c <= 9'b101011111;
				8'b1101000: c <= 9'b110110;
				8'b101100: c <= 9'b11000111;
				8'b100100: c <= 9'b101001;
				8'b1111000: c <= 9'b111001010;
				8'b1000101: c <= 9'b1100110;
				8'b1011001: c <= 9'b11110101;
				8'b110100: c <= 9'b101010;
				8'b1111001: c <= 9'b101100;
				8'b1110001: c <= 9'b1011110;
				8'b1001111: c <= 9'b111101001;
				8'b1100101: c <= 9'b111011100;
				8'b1111110: c <= 9'b11101000;
				8'b1111100: c <= 9'b100001001;
				8'b1010110: c <= 9'b11001001;
				8'b110010: c <= 9'b110010101;
				8'b1101101: c <= 9'b101011000;
				8'b100011: c <= 9'b101101;
				8'b1110101: c <= 9'b1000111;
				8'b1111101: c <= 9'b110011;
				8'b101001: c <= 9'b1011010;
				8'b1010010: c <= 9'b110011;
				8'b1011000: c <= 9'b101111001;
				8'b101110: c <= 9'b101001000;
				8'b1000001: c <= 9'b111000110;
				default: c <= 9'b0;
			endcase
			9'b1100010 : case(di)
				8'b1000011: c <= 9'b101010010;
				8'b101000: c <= 9'b1001;
				8'b111010: c <= 9'b101010;
				8'b110110: c <= 9'b10100;
				8'b1100100: c <= 9'b111101001;
				8'b1000000: c <= 9'b11011010;
				8'b1110110: c <= 9'b111100100;
				8'b100101: c <= 9'b111110110;
				8'b101111: c <= 9'b100010101;
				8'b100110: c <= 9'b11010011;
				8'b1100011: c <= 9'b10111101;
				8'b1001000: c <= 9'b100011100;
				8'b111000: c <= 9'b111001001;
				8'b110001: c <= 9'b11101101;
				8'b1010111: c <= 9'b1100001;
				8'b1001110: c <= 9'b100110010;
				8'b1101010: c <= 9'b110100010;
				8'b1001001: c <= 9'b101100011;
				8'b1100000: c <= 9'b1111100;
				8'b110111: c <= 9'b10110111;
				8'b1011101: c <= 9'b11011;
				8'b1011011: c <= 9'b111111000;
				8'b111001: c <= 9'b110110;
				8'b1001010: c <= 9'b110010111;
				8'b110011: c <= 9'b111101110;
				8'b1101100: c <= 9'b11001011;
				8'b1110111: c <= 9'b111001;
				8'b101011: c <= 9'b111000011;
				8'b1101011: c <= 9'b100101000;
				8'b111100: c <= 9'b110011101;
				8'b1000111: c <= 9'b111100110;
				8'b1011111: c <= 9'b111100001;
				8'b1110100: c <= 9'b10101010;
				8'b101101: c <= 9'b10011001;
				8'b1010011: c <= 9'b111000110;
				8'b1100001: c <= 9'b1001100;
				8'b110101: c <= 9'b11100101;
				8'b1000100: c <= 9'b110011011;
				8'b1010001: c <= 9'b11001100;
				8'b1010100: c <= 9'b1101111;
				8'b1100110: c <= 9'b110000110;
				8'b101010: c <= 9'b100001100;
				8'b1011110: c <= 9'b11111001;
				8'b1100111: c <= 9'b11000111;
				8'b1011010: c <= 9'b1010010;
				8'b1000010: c <= 9'b100101000;
				8'b111101: c <= 9'b11000001;
				8'b110000: c <= 9'b10010111;
				8'b111110: c <= 9'b100110111;
				8'b1100010: c <= 9'b110001110;
				8'b1110000: c <= 9'b100100101;
				8'b1101001: c <= 9'b100001010;
				8'b1110011: c <= 9'b10111011;
				8'b1001100: c <= 9'b111100011;
				8'b100001: c <= 9'b1101000;
				8'b1000110: c <= 9'b1001110;
				8'b1110010: c <= 9'b11110001;
				8'b1010000: c <= 9'b1111110;
				8'b1111010: c <= 9'b11010101;
				8'b1010101: c <= 9'b110111000;
				8'b111011: c <= 9'b10110101;
				8'b1001101: c <= 9'b11111;
				8'b111111: c <= 9'b100011111;
				8'b1101110: c <= 9'b100001110;
				8'b1111011: c <= 9'b101110101;
				8'b1001011: c <= 9'b100100011;
				8'b1101111: c <= 9'b1101101;
				8'b1101000: c <= 9'b1001010;
				8'b101100: c <= 9'b11010100;
				8'b100100: c <= 9'b10111010;
				8'b1111000: c <= 9'b11000110;
				8'b1000101: c <= 9'b10110;
				8'b1011001: c <= 9'b111010111;
				8'b110100: c <= 9'b101010000;
				8'b1111001: c <= 9'b100001101;
				8'b1110001: c <= 9'b100010111;
				8'b1001111: c <= 9'b101110;
				8'b1100101: c <= 9'b100011111;
				8'b1111110: c <= 9'b11101000;
				8'b1111100: c <= 9'b111011001;
				8'b1010110: c <= 9'b110111011;
				8'b110010: c <= 9'b1010101;
				8'b1101101: c <= 9'b10101110;
				8'b100011: c <= 9'b101101110;
				8'b1110101: c <= 9'b1101110;
				8'b1111101: c <= 9'b111100000;
				8'b101001: c <= 9'b11101;
				8'b1010010: c <= 9'b1010101;
				8'b1011000: c <= 9'b111100101;
				8'b101110: c <= 9'b1100101;
				8'b1000001: c <= 9'b11101100;
				default: c <= 9'b0;
			endcase
			9'b1110111 : case(di)
				8'b1000011: c <= 9'b111011;
				8'b101000: c <= 9'b1100001;
				8'b111010: c <= 9'b1111;
				8'b110110: c <= 9'b1001101;
				8'b1100100: c <= 9'b11111;
				8'b1000000: c <= 9'b11010100;
				8'b1110110: c <= 9'b101000001;
				8'b100101: c <= 9'b10100000;
				8'b101111: c <= 9'b10010001;
				8'b100110: c <= 9'b100101110;
				8'b1100011: c <= 9'b101111111;
				8'b1001000: c <= 9'b100101010;
				8'b111000: c <= 9'b100111010;
				8'b110001: c <= 9'b10101110;
				8'b1010111: c <= 9'b101100111;
				8'b1001110: c <= 9'b111100010;
				8'b1101010: c <= 9'b110001010;
				8'b1001001: c <= 9'b101001011;
				8'b1100000: c <= 9'b10101011;
				8'b110111: c <= 9'b11010111;
				8'b1011101: c <= 9'b111110000;
				8'b1011011: c <= 9'b100011100;
				8'b111001: c <= 9'b1010010;
				8'b1001010: c <= 9'b1001110;
				8'b110011: c <= 9'b1100000;
				8'b1101100: c <= 9'b111101001;
				8'b1110111: c <= 9'b111011011;
				8'b101011: c <= 9'b100010;
				8'b1101011: c <= 9'b10110001;
				8'b111100: c <= 9'b11101001;
				8'b1000111: c <= 9'b111100001;
				8'b1011111: c <= 9'b110000101;
				8'b1110100: c <= 9'b110110011;
				8'b101101: c <= 9'b11111010;
				8'b1010011: c <= 9'b11110;
				8'b1100001: c <= 9'b100110111;
				8'b110101: c <= 9'b111101111;
				8'b1000100: c <= 9'b1010000;
				8'b1010001: c <= 9'b1110010;
				8'b1010100: c <= 9'b111010100;
				8'b1100110: c <= 9'b10101000;
				8'b101010: c <= 9'b101010011;
				8'b1011110: c <= 9'b110111110;
				8'b1100111: c <= 9'b10000101;
				8'b1011010: c <= 9'b10;
				8'b1000010: c <= 9'b111000;
				8'b111101: c <= 9'b101000010;
				8'b110000: c <= 9'b111011110;
				8'b111110: c <= 9'b101010010;
				8'b1100010: c <= 9'b101110110;
				8'b1110000: c <= 9'b10001000;
				8'b1101001: c <= 9'b111001010;
				8'b1110011: c <= 9'b10110;
				8'b1001100: c <= 9'b100011000;
				8'b100001: c <= 9'b1010001;
				8'b1000110: c <= 9'b111001001;
				8'b1110010: c <= 9'b110011110;
				8'b1010000: c <= 9'b11101000;
				8'b1111010: c <= 9'b100100000;
				8'b1010101: c <= 9'b10011100;
				8'b111011: c <= 9'b10100000;
				8'b1001101: c <= 9'b110100110;
				8'b111111: c <= 9'b100010110;
				8'b1101110: c <= 9'b101001111;
				8'b1111011: c <= 9'b1110011;
				8'b1001011: c <= 9'b110101011;
				8'b1101111: c <= 9'b110110111;
				8'b1101000: c <= 9'b10000;
				8'b101100: c <= 9'b1010011;
				8'b100100: c <= 9'b10011;
				8'b1111000: c <= 9'b110100111;
				8'b1000101: c <= 9'b111111010;
				8'b1011001: c <= 9'b10010001;
				8'b110100: c <= 9'b110101;
				8'b1111001: c <= 9'b101000010;
				8'b1110001: c <= 9'b100010100;
				8'b1001111: c <= 9'b11011011;
				8'b1100101: c <= 9'b10;
				8'b1111110: c <= 9'b100111010;
				8'b1111100: c <= 9'b1111;
				8'b1010110: c <= 9'b100111;
				8'b110010: c <= 9'b100011010;
				8'b1101101: c <= 9'b100;
				8'b100011: c <= 9'b10010011;
				8'b1110101: c <= 9'b101110100;
				8'b1111101: c <= 9'b111001010;
				8'b101001: c <= 9'b100001111;
				8'b1010010: c <= 9'b110101;
				8'b1011000: c <= 9'b10110110;
				8'b101110: c <= 9'b111000111;
				8'b1000001: c <= 9'b110000001;
				default: c <= 9'b0;
			endcase
			9'b1111 : case(di)
				8'b1000011: c <= 9'b101100110;
				8'b101000: c <= 9'b11010101;
				8'b111010: c <= 9'b10100010;
				8'b110110: c <= 9'b110010010;
				8'b1100100: c <= 9'b111000111;
				8'b1000000: c <= 9'b1100110;
				8'b1110110: c <= 9'b101001001;
				8'b100101: c <= 9'b101000101;
				8'b101111: c <= 9'b101011001;
				8'b100110: c <= 9'b10001111;
				8'b1100011: c <= 9'b10010011;
				8'b1001000: c <= 9'b1110101;
				8'b111000: c <= 9'b100001101;
				8'b110001: c <= 9'b111000;
				8'b1010111: c <= 9'b111100;
				8'b1001110: c <= 9'b100111110;
				8'b1101010: c <= 9'b10111111;
				8'b1001001: c <= 9'b101000111;
				8'b1100000: c <= 9'b111001011;
				8'b110111: c <= 9'b1111100;
				8'b1011101: c <= 9'b111110011;
				8'b1011011: c <= 9'b100000111;
				8'b111001: c <= 9'b110100101;
				8'b1001010: c <= 9'b10101111;
				8'b110011: c <= 9'b10111111;
				8'b1101100: c <= 9'b111010000;
				8'b1110111: c <= 9'b11010001;
				8'b101011: c <= 9'b111001101;
				8'b1101011: c <= 9'b111111000;
				8'b111100: c <= 9'b101111010;
				8'b1000111: c <= 9'b110001110;
				8'b1011111: c <= 9'b111000100;
				8'b1110100: c <= 9'b100000110;
				8'b101101: c <= 9'b100001110;
				8'b1010011: c <= 9'b10011001;
				8'b1100001: c <= 9'b1110000;
				8'b110101: c <= 9'b11111;
				8'b1000100: c <= 9'b111111010;
				8'b1010001: c <= 9'b100100000;
				8'b1010100: c <= 9'b100101001;
				8'b1100110: c <= 9'b101100100;
				8'b101010: c <= 9'b100000011;
				8'b1011110: c <= 9'b101000100;
				8'b1100111: c <= 9'b11000100;
				8'b1011010: c <= 9'b110100100;
				8'b1000010: c <= 9'b11111;
				8'b111101: c <= 9'b111011001;
				8'b110000: c <= 9'b10100100;
				8'b111110: c <= 9'b110100101;
				8'b1100010: c <= 9'b111111101;
				8'b1110000: c <= 9'b1111100;
				8'b1101001: c <= 9'b11100010;
				8'b1110011: c <= 9'b11011011;
				8'b1001100: c <= 9'b10110010;
				8'b100001: c <= 9'b100111;
				8'b1000110: c <= 9'b110000110;
				8'b1110010: c <= 9'b111111101;
				8'b1010000: c <= 9'b111010000;
				8'b1111010: c <= 9'b111110101;
				8'b1010101: c <= 9'b11100101;
				8'b111011: c <= 9'b100000000;
				8'b1001101: c <= 9'b11111110;
				8'b111111: c <= 9'b101101000;
				8'b1101110: c <= 9'b111101101;
				8'b1111011: c <= 9'b11000111;
				8'b1001011: c <= 9'b110100111;
				8'b1101111: c <= 9'b111100100;
				8'b1101000: c <= 9'b1010000;
				8'b101100: c <= 9'b11100111;
				8'b100100: c <= 9'b101000101;
				8'b1111000: c <= 9'b10010110;
				8'b1000101: c <= 9'b101010110;
				8'b1011001: c <= 9'b101101000;
				8'b110100: c <= 9'b11011101;
				8'b1111001: c <= 9'b110110100;
				8'b1110001: c <= 9'b110110110;
				8'b1001111: c <= 9'b111100001;
				8'b1100101: c <= 9'b111101;
				8'b1111110: c <= 9'b110011011;
				8'b1111100: c <= 9'b100011000;
				8'b1010110: c <= 9'b101100001;
				8'b110010: c <= 9'b111111001;
				8'b1101101: c <= 9'b101001110;
				8'b100011: c <= 9'b101101101;
				8'b1110101: c <= 9'b111000111;
				8'b1111101: c <= 9'b11000011;
				8'b101001: c <= 9'b10100010;
				8'b1010010: c <= 9'b100001001;
				8'b1011000: c <= 9'b100011100;
				8'b101110: c <= 9'b10000110;
				8'b1000001: c <= 9'b110100110;
				default: c <= 9'b0;
			endcase
			9'b11100111 : case(di)
				8'b1000011: c <= 9'b111001011;
				8'b101000: c <= 9'b101000;
				8'b111010: c <= 9'b101100;
				8'b110110: c <= 9'b101111001;
				8'b1100100: c <= 9'b100111100;
				8'b1000000: c <= 9'b10011;
				8'b1110110: c <= 9'b101101111;
				8'b100101: c <= 9'b1111010;
				8'b101111: c <= 9'b1101000;
				8'b100110: c <= 9'b101010111;
				8'b1100011: c <= 9'b1111011;
				8'b1001000: c <= 9'b110100001;
				8'b111000: c <= 9'b1001011;
				8'b110001: c <= 9'b11110101;
				8'b1010111: c <= 9'b111111111;
				8'b1001110: c <= 9'b100000011;
				8'b1101010: c <= 9'b11100001;
				8'b1001001: c <= 9'b10111;
				8'b1100000: c <= 9'b10111110;
				8'b110111: c <= 9'b1111010;
				8'b1011101: c <= 9'b11011110;
				8'b1011011: c <= 9'b11000100;
				8'b111001: c <= 9'b111001100;
				8'b1001010: c <= 9'b10111010;
				8'b110011: c <= 9'b1100100;
				8'b1101100: c <= 9'b11010;
				8'b1110111: c <= 9'b10001100;
				8'b101011: c <= 9'b10111010;
				8'b1101011: c <= 9'b1011010;
				8'b111100: c <= 9'b11101;
				8'b1000111: c <= 9'b11101011;
				8'b1011111: c <= 9'b100010010;
				8'b1110100: c <= 9'b111110011;
				8'b101101: c <= 9'b100001010;
				8'b1010011: c <= 9'b100101100;
				8'b1100001: c <= 9'b110010110;
				8'b110101: c <= 9'b10001111;
				8'b1000100: c <= 9'b101101111;
				8'b1010001: c <= 9'b111101100;
				8'b1010100: c <= 9'b10101000;
				8'b1100110: c <= 9'b111000101;
				8'b101010: c <= 9'b1100110;
				8'b1011110: c <= 9'b111100100;
				8'b1100111: c <= 9'b101101100;
				8'b1011010: c <= 9'b110001;
				8'b1000010: c <= 9'b1111111;
				8'b111101: c <= 9'b10011001;
				8'b110000: c <= 9'b11111100;
				8'b111110: c <= 9'b110011110;
				8'b1100010: c <= 9'b1011111;
				8'b1110000: c <= 9'b101111110;
				8'b1101001: c <= 9'b110010101;
				8'b1110011: c <= 9'b100111010;
				8'b1001100: c <= 9'b10001101;
				8'b100001: c <= 9'b10001000;
				8'b1000110: c <= 9'b10111110;
				8'b1110010: c <= 9'b101100011;
				8'b1010000: c <= 9'b110011111;
				8'b1111010: c <= 9'b1000010;
				8'b1010101: c <= 9'b110011010;
				8'b111011: c <= 9'b111101110;
				8'b1001101: c <= 9'b101011110;
				8'b111111: c <= 9'b101000;
				8'b1101110: c <= 9'b111001001;
				8'b1111011: c <= 9'b10;
				8'b1001011: c <= 9'b110111010;
				8'b1101111: c <= 9'b111011101;
				8'b1101000: c <= 9'b11101000;
				8'b101100: c <= 9'b110011011;
				8'b100100: c <= 9'b1100011;
				8'b1111000: c <= 9'b100111111;
				8'b1000101: c <= 9'b10001001;
				8'b1011001: c <= 9'b101100010;
				8'b110100: c <= 9'b10101;
				8'b1111001: c <= 9'b101100011;
				8'b1110001: c <= 9'b1000100;
				8'b1001111: c <= 9'b11000100;
				8'b1100101: c <= 9'b1100101;
				8'b1111110: c <= 9'b101001011;
				8'b1111100: c <= 9'b100110011;
				8'b1010110: c <= 9'b101110101;
				8'b110010: c <= 9'b111111111;
				8'b1101101: c <= 9'b11100110;
				8'b100011: c <= 9'b1001001;
				8'b1110101: c <= 9'b11100;
				8'b1111101: c <= 9'b111100100;
				8'b101001: c <= 9'b1110111;
				8'b1010010: c <= 9'b10001000;
				8'b1011000: c <= 9'b10111011;
				8'b101110: c <= 9'b110111011;
				8'b1000001: c <= 9'b101110110;
				default: c <= 9'b0;
			endcase
			9'b1100 : case(di)
				8'b1000011: c <= 9'b1110100;
				8'b101000: c <= 9'b100000010;
				8'b111010: c <= 9'b111111010;
				8'b110110: c <= 9'b100110101;
				8'b1100100: c <= 9'b1110011;
				8'b1000000: c <= 9'b110100100;
				8'b1110110: c <= 9'b101011110;
				8'b100101: c <= 9'b101011000;
				8'b101111: c <= 9'b11011001;
				8'b100110: c <= 9'b100001;
				8'b1100011: c <= 9'b110111000;
				8'b1001000: c <= 9'b110011101;
				8'b111000: c <= 9'b100010000;
				8'b110001: c <= 9'b1010111;
				8'b1010111: c <= 9'b11111110;
				8'b1001110: c <= 9'b110101110;
				8'b1101010: c <= 9'b100000000;
				8'b1001001: c <= 9'b110101111;
				8'b1100000: c <= 9'b100101001;
				8'b110111: c <= 9'b101010110;
				8'b1011101: c <= 9'b111101111;
				8'b1011011: c <= 9'b1011000;
				8'b111001: c <= 9'b10011001;
				8'b1001010: c <= 9'b1110111;
				8'b110011: c <= 9'b1011011;
				8'b1101100: c <= 9'b111001011;
				8'b1110111: c <= 9'b111101000;
				8'b101011: c <= 9'b1110;
				8'b1101011: c <= 9'b10111111;
				8'b111100: c <= 9'b1000101;
				8'b1000111: c <= 9'b101011;
				8'b1011111: c <= 9'b10111100;
				8'b1110100: c <= 9'b1011100;
				8'b101101: c <= 9'b10101110;
				8'b1010011: c <= 9'b10110011;
				8'b1100001: c <= 9'b11010000;
				8'b110101: c <= 9'b1101101;
				8'b1000100: c <= 9'b101000100;
				8'b1010001: c <= 9'b111000100;
				8'b1010100: c <= 9'b100101101;
				8'b1100110: c <= 9'b10001011;
				8'b101010: c <= 9'b101110101;
				8'b1011110: c <= 9'b111001110;
				8'b1100111: c <= 9'b110010101;
				8'b1011010: c <= 9'b11011100;
				8'b1000010: c <= 9'b10010000;
				8'b111101: c <= 9'b101100100;
				8'b110000: c <= 9'b11110001;
				8'b111110: c <= 9'b1111000;
				8'b1100010: c <= 9'b101010100;
				8'b1110000: c <= 9'b100000011;
				8'b1101001: c <= 9'b11001000;
				8'b1110011: c <= 9'b10110010;
				8'b1001100: c <= 9'b100100;
				8'b100001: c <= 9'b101110000;
				8'b1000110: c <= 9'b11111010;
				8'b1110010: c <= 9'b100001;
				8'b1010000: c <= 9'b111001101;
				8'b1111010: c <= 9'b110001001;
				8'b1010101: c <= 9'b1101100;
				8'b111011: c <= 9'b111100101;
				8'b1001101: c <= 9'b101111111;
				8'b111111: c <= 9'b111000;
				8'b1101110: c <= 9'b1111010;
				8'b1111011: c <= 9'b11111010;
				8'b1001011: c <= 9'b100110111;
				8'b1101111: c <= 9'b100101011;
				8'b1101000: c <= 9'b11111011;
				8'b101100: c <= 9'b100111100;
				8'b100100: c <= 9'b110010010;
				8'b1111000: c <= 9'b11100111;
				8'b1000101: c <= 9'b110010110;
				8'b1011001: c <= 9'b100101000;
				8'b110100: c <= 9'b100010111;
				8'b1111001: c <= 9'b110010;
				8'b1110001: c <= 9'b11100011;
				8'b1001111: c <= 9'b111000101;
				8'b1100101: c <= 9'b11011000;
				8'b1111110: c <= 9'b110001000;
				8'b1111100: c <= 9'b101101010;
				8'b1010110: c <= 9'b10010;
				8'b110010: c <= 9'b110101111;
				8'b1101101: c <= 9'b11001110;
				8'b100011: c <= 9'b110010100;
				8'b1110101: c <= 9'b100001;
				8'b1111101: c <= 9'b10010101;
				8'b101001: c <= 9'b100101101;
				8'b1010010: c <= 9'b111001110;
				8'b1011000: c <= 9'b10000011;
				8'b101110: c <= 9'b10110;
				8'b1000001: c <= 9'b111011101;
				default: c <= 9'b0;
			endcase
			9'b11011001 : case(di)
				8'b1000011: c <= 9'b1010011;
				8'b101000: c <= 9'b111101111;
				8'b111010: c <= 9'b101011110;
				8'b110110: c <= 9'b101100001;
				8'b1100100: c <= 9'b10111001;
				8'b1000000: c <= 9'b11111;
				8'b1110110: c <= 9'b101000101;
				8'b100101: c <= 9'b111001010;
				8'b101111: c <= 9'b11000111;
				8'b100110: c <= 9'b11100011;
				8'b1100011: c <= 9'b101000100;
				8'b1001000: c <= 9'b10000101;
				8'b111000: c <= 9'b1101001;
				8'b110001: c <= 9'b110001001;
				8'b1010111: c <= 9'b1110001;
				8'b1001110: c <= 9'b110011001;
				8'b1101010: c <= 9'b11110110;
				8'b1001001: c <= 9'b100011000;
				8'b1100000: c <= 9'b110100010;
				8'b110111: c <= 9'b101011010;
				8'b1011101: c <= 9'b11110011;
				8'b1011011: c <= 9'b110001101;
				8'b111001: c <= 9'b11011011;
				8'b1001010: c <= 9'b100000000;
				8'b110011: c <= 9'b110000;
				8'b1101100: c <= 9'b101010010;
				8'b1110111: c <= 9'b10011101;
				8'b101011: c <= 9'b110001110;
				8'b1101011: c <= 9'b100;
				8'b111100: c <= 9'b101001111;
				8'b1000111: c <= 9'b110111100;
				8'b1011111: c <= 9'b10011111;
				8'b1110100: c <= 9'b1011111;
				8'b101101: c <= 9'b110100011;
				8'b1010011: c <= 9'b10101000;
				8'b1100001: c <= 9'b10111010;
				8'b110101: c <= 9'b10001111;
				8'b1000100: c <= 9'b1100100;
				8'b1010001: c <= 9'b11101011;
				8'b1010100: c <= 9'b101000110;
				8'b1100110: c <= 9'b1100000;
				8'b101010: c <= 9'b101000110;
				8'b1011110: c <= 9'b111101110;
				8'b1100111: c <= 9'b101010010;
				8'b1011010: c <= 9'b101100101;
				8'b1000010: c <= 9'b110110011;
				8'b111101: c <= 9'b101101100;
				8'b110000: c <= 9'b1001;
				8'b111110: c <= 9'b1111001;
				8'b1100010: c <= 9'b101100100;
				8'b1110000: c <= 9'b10100101;
				8'b1101001: c <= 9'b100100010;
				8'b1110011: c <= 9'b110111110;
				8'b1001100: c <= 9'b1110101;
				8'b100001: c <= 9'b110110101;
				8'b1000110: c <= 9'b101001111;
				8'b1110010: c <= 9'b1101111;
				8'b1010000: c <= 9'b100010010;
				8'b1111010: c <= 9'b110000101;
				8'b1010101: c <= 9'b10110010;
				8'b111011: c <= 9'b110010010;
				8'b1001101: c <= 9'b111111010;
				8'b111111: c <= 9'b1101110;
				8'b1101110: c <= 9'b100100010;
				8'b1111011: c <= 9'b10000110;
				8'b1001011: c <= 9'b111101111;
				8'b1101111: c <= 9'b1111010;
				8'b1101000: c <= 9'b101100000;
				8'b101100: c <= 9'b110000110;
				8'b100100: c <= 9'b11101001;
				8'b1111000: c <= 9'b110110100;
				8'b1000101: c <= 9'b111010110;
				8'b1011001: c <= 9'b11011100;
				8'b110100: c <= 9'b11001100;
				8'b1111001: c <= 9'b101010101;
				8'b1110001: c <= 9'b110101;
				8'b1001111: c <= 9'b111011001;
				8'b1100101: c <= 9'b10100010;
				8'b1111110: c <= 9'b110110011;
				8'b1111100: c <= 9'b101101100;
				8'b1010110: c <= 9'b10010;
				8'b110010: c <= 9'b110100001;
				8'b1101101: c <= 9'b111011001;
				8'b100011: c <= 9'b110101001;
				8'b1110101: c <= 9'b101101000;
				8'b1111101: c <= 9'b100101011;
				8'b101001: c <= 9'b111100100;
				8'b1010010: c <= 9'b1000001;
				8'b1011000: c <= 9'b11011101;
				8'b101110: c <= 9'b11010101;
				8'b1000001: c <= 9'b10111;
				default: c <= 9'b0;
			endcase
			9'b10111111 : case(di)
				8'b1000011: c <= 9'b11101001;
				8'b101000: c <= 9'b100000100;
				8'b111010: c <= 9'b101111000;
				8'b110110: c <= 9'b110101111;
				8'b1100100: c <= 9'b111001001;
				8'b1000000: c <= 9'b10000;
				8'b1110110: c <= 9'b111000101;
				8'b100101: c <= 9'b10010110;
				8'b101111: c <= 9'b10000111;
				8'b100110: c <= 9'b111000011;
				8'b1100011: c <= 9'b110;
				8'b1001000: c <= 9'b10011000;
				8'b111000: c <= 9'b10101110;
				8'b110001: c <= 9'b110011111;
				8'b1010111: c <= 9'b10100111;
				8'b1001110: c <= 9'b10111001;
				8'b1101010: c <= 9'b100001101;
				8'b1001001: c <= 9'b111100;
				8'b1100000: c <= 9'b1111000;
				8'b110111: c <= 9'b100101110;
				8'b1011101: c <= 9'b10001101;
				8'b1011011: c <= 9'b100010;
				8'b111001: c <= 9'b100001111;
				8'b1001010: c <= 9'b100100000;
				8'b110011: c <= 9'b100100010;
				8'b1101100: c <= 9'b110110010;
				8'b1110111: c <= 9'b110001000;
				8'b101011: c <= 9'b110001001;
				8'b1101011: c <= 9'b110011001;
				8'b111100: c <= 9'b10011111;
				8'b1000111: c <= 9'b101010110;
				8'b1011111: c <= 9'b10011011;
				8'b1110100: c <= 9'b1110001;
				8'b101101: c <= 9'b11110;
				8'b1010011: c <= 9'b101010000;
				8'b1100001: c <= 9'b1010001;
				8'b110101: c <= 9'b110111001;
				8'b1000100: c <= 9'b1101000;
				8'b1010001: c <= 9'b11101;
				8'b1010100: c <= 9'b10010111;
				8'b1100110: c <= 9'b110100110;
				8'b101010: c <= 9'b11;
				8'b1011110: c <= 9'b111011111;
				8'b1100111: c <= 9'b1101100;
				8'b1011010: c <= 9'b111010010;
				8'b1000010: c <= 9'b10001111;
				8'b111101: c <= 9'b11101001;
				8'b110000: c <= 9'b1111101;
				8'b111110: c <= 9'b101101010;
				8'b1100010: c <= 9'b111001000;
				8'b1110000: c <= 9'b100001;
				8'b1101001: c <= 9'b100110100;
				8'b1110011: c <= 9'b110100000;
				8'b1001100: c <= 9'b111101101;
				8'b100001: c <= 9'b100111111;
				8'b1000110: c <= 9'b1110011;
				8'b1110010: c <= 9'b100110011;
				8'b1010000: c <= 9'b111010001;
				8'b1111010: c <= 9'b100011111;
				8'b1010101: c <= 9'b11011100;
				8'b111011: c <= 9'b111011111;
				8'b1001101: c <= 9'b111000100;
				8'b111111: c <= 9'b110010110;
				8'b1101110: c <= 9'b101100001;
				8'b1111011: c <= 9'b1100110;
				8'b1001011: c <= 9'b10011010;
				8'b1101111: c <= 9'b110001;
				8'b1101000: c <= 9'b10110011;
				8'b101100: c <= 9'b100111100;
				8'b100100: c <= 9'b10001001;
				8'b1111000: c <= 9'b111011110;
				8'b1000101: c <= 9'b11001111;
				8'b1011001: c <= 9'b111100010;
				8'b110100: c <= 9'b100110;
				8'b1111001: c <= 9'b11101001;
				8'b1110001: c <= 9'b101110001;
				8'b1001111: c <= 9'b110010100;
				8'b1100101: c <= 9'b10111101;
				8'b1111110: c <= 9'b11011001;
				8'b1111100: c <= 9'b100111101;
				8'b1010110: c <= 9'b11100010;
				8'b110010: c <= 9'b11;
				8'b1101101: c <= 9'b10100101;
				8'b100011: c <= 9'b101010001;
				8'b1110101: c <= 9'b11001101;
				8'b1111101: c <= 9'b11101100;
				8'b101001: c <= 9'b111001011;
				8'b1010010: c <= 9'b100111000;
				8'b1011000: c <= 9'b110011110;
				8'b101110: c <= 9'b111011110;
				8'b1000001: c <= 9'b101110101;
				default: c <= 9'b0;
			endcase
			9'b101010110 : case(di)
				8'b1000011: c <= 9'b111101110;
				8'b101000: c <= 9'b10101001;
				8'b111010: c <= 9'b100110;
				8'b110110: c <= 9'b111010100;
				8'b1100100: c <= 9'b111000100;
				8'b1000000: c <= 9'b11010001;
				8'b1110110: c <= 9'b10101011;
				8'b100101: c <= 9'b11100011;
				8'b101111: c <= 9'b100101001;
				8'b100110: c <= 9'b11100110;
				8'b1100011: c <= 9'b1011011;
				8'b1001000: c <= 9'b110001000;
				8'b111000: c <= 9'b10001111;
				8'b110001: c <= 9'b110101101;
				8'b1010111: c <= 9'b111101100;
				8'b1001110: c <= 9'b100001010;
				8'b1101010: c <= 9'b101111110;
				8'b1001001: c <= 9'b111000010;
				8'b1100000: c <= 9'b1101001;
				8'b110111: c <= 9'b100111100;
				8'b1011101: c <= 9'b11100;
				8'b1011011: c <= 9'b1001000;
				8'b111001: c <= 9'b101101100;
				8'b1001010: c <= 9'b100011101;
				8'b110011: c <= 9'b11001100;
				8'b1101100: c <= 9'b110111001;
				8'b1110111: c <= 9'b10010100;
				8'b101011: c <= 9'b10011;
				8'b1101011: c <= 9'b110011010;
				8'b111100: c <= 9'b10000;
				8'b1000111: c <= 9'b1010001;
				8'b1011111: c <= 9'b10101010;
				8'b1110100: c <= 9'b1100011;
				8'b101101: c <= 9'b111101110;
				8'b1010011: c <= 9'b100010010;
				8'b1100001: c <= 9'b100101001;
				8'b110101: c <= 9'b11101100;
				8'b1000100: c <= 9'b10110010;
				8'b1010001: c <= 9'b111111111;
				8'b1010100: c <= 9'b111100101;
				8'b1100110: c <= 9'b111000110;
				8'b101010: c <= 9'b1110111;
				8'b1011110: c <= 9'b101111010;
				8'b1100111: c <= 9'b11001001;
				8'b1011010: c <= 9'b111111000;
				8'b1000010: c <= 9'b110111001;
				8'b111101: c <= 9'b111001110;
				8'b110000: c <= 9'b110110011;
				8'b111110: c <= 9'b101011010;
				8'b1100010: c <= 9'b111101;
				8'b1110000: c <= 9'b1111001;
				8'b1101001: c <= 9'b111111001;
				8'b1110011: c <= 9'b101111111;
				8'b1001100: c <= 9'b11110010;
				8'b100001: c <= 9'b111110000;
				8'b1000110: c <= 9'b110001001;
				8'b1110010: c <= 9'b101111001;
				8'b1010000: c <= 9'b111000000;
				8'b1111010: c <= 9'b110110000;
				8'b1010101: c <= 9'b11101100;
				8'b111011: c <= 9'b10010111;
				8'b1001101: c <= 9'b111011010;
				8'b111111: c <= 9'b110000111;
				8'b1101110: c <= 9'b100101010;
				8'b1111011: c <= 9'b1011100;
				8'b1001011: c <= 9'b110010111;
				8'b1101111: c <= 9'b101010011;
				8'b1101000: c <= 9'b100010101;
				8'b101100: c <= 9'b101000;
				8'b100100: c <= 9'b1000;
				8'b1111000: c <= 9'b11010100;
				8'b1000101: c <= 9'b11011;
				8'b1011001: c <= 9'b110100101;
				8'b110100: c <= 9'b10000111;
				8'b1111001: c <= 9'b100000100;
				8'b1110001: c <= 9'b111010111;
				8'b1001111: c <= 9'b1010101;
				8'b1100101: c <= 9'b111000000;
				8'b1111110: c <= 9'b1101000;
				8'b1111100: c <= 9'b100101010;
				8'b1010110: c <= 9'b111000010;
				8'b110010: c <= 9'b11011001;
				8'b1101101: c <= 9'b101001010;
				8'b100011: c <= 9'b100100001;
				8'b1110101: c <= 9'b100010101;
				8'b1111101: c <= 9'b1000101;
				8'b101001: c <= 9'b100000101;
				8'b1010010: c <= 9'b101010101;
				8'b1011000: c <= 9'b11111000;
				8'b101110: c <= 9'b11111100;
				8'b1000001: c <= 9'b10101111;
				default: c <= 9'b0;
			endcase
			9'b10011100 : case(di)
				8'b1000011: c <= 9'b100011011;
				8'b101000: c <= 9'b101011001;
				8'b111010: c <= 9'b10010011;
				8'b110110: c <= 9'b101100010;
				8'b1100100: c <= 9'b10110110;
				8'b1000000: c <= 9'b101101001;
				8'b1110110: c <= 9'b10110100;
				8'b100101: c <= 9'b1000001;
				8'b101111: c <= 9'b10111100;
				8'b100110: c <= 9'b101100000;
				8'b1100011: c <= 9'b10010110;
				8'b1001000: c <= 9'b1010000;
				8'b111000: c <= 9'b100101000;
				8'b110001: c <= 9'b100101;
				8'b1010111: c <= 9'b101110111;
				8'b1001110: c <= 9'b10001111;
				8'b1101010: c <= 9'b100001;
				8'b1001001: c <= 9'b101010110;
				8'b1100000: c <= 9'b111001111;
				8'b110111: c <= 9'b100101011;
				8'b1011101: c <= 9'b101010011;
				8'b1011011: c <= 9'b110101110;
				8'b111001: c <= 9'b101000001;
				8'b1001010: c <= 9'b110101111;
				8'b110011: c <= 9'b111110101;
				8'b1101100: c <= 9'b100101101;
				8'b1110111: c <= 9'b10111000;
				8'b101011: c <= 9'b10010000;
				8'b1101011: c <= 9'b101101111;
				8'b111100: c <= 9'b101100101;
				8'b1000111: c <= 9'b11100100;
				8'b1011111: c <= 9'b11110100;
				8'b1110100: c <= 9'b10;
				8'b101101: c <= 9'b100101110;
				8'b1010011: c <= 9'b10000111;
				8'b1100001: c <= 9'b10110011;
				8'b110101: c <= 9'b101100001;
				8'b1000100: c <= 9'b101010110;
				8'b1010001: c <= 9'b111001100;
				8'b1010100: c <= 9'b11101100;
				8'b1100110: c <= 9'b11011110;
				8'b101010: c <= 9'b110010100;
				8'b1011110: c <= 9'b11100110;
				8'b1100111: c <= 9'b100001;
				8'b1011010: c <= 9'b11010001;
				8'b1000010: c <= 9'b10101001;
				8'b111101: c <= 9'b111100001;
				8'b110000: c <= 9'b100001010;
				8'b111110: c <= 9'b101011011;
				8'b1100010: c <= 9'b100000110;
				8'b1110000: c <= 9'b1000011;
				8'b1101001: c <= 9'b1110011;
				8'b1110011: c <= 9'b1100011;
				8'b1001100: c <= 9'b100010001;
				8'b100001: c <= 9'b100110101;
				8'b1000110: c <= 9'b11010010;
				8'b1110010: c <= 9'b100001101;
				8'b1010000: c <= 9'b110111111;
				8'b1111010: c <= 9'b110010011;
				8'b1010101: c <= 9'b110101001;
				8'b111011: c <= 9'b100001011;
				8'b1001101: c <= 9'b1100001;
				8'b111111: c <= 9'b111110000;
				8'b1101110: c <= 9'b11111011;
				8'b1111011: c <= 9'b11000000;
				8'b1001011: c <= 9'b101110000;
				8'b1101111: c <= 9'b101100101;
				8'b1101000: c <= 9'b101010011;
				8'b101100: c <= 9'b111011011;
				8'b100100: c <= 9'b110100010;
				8'b1111000: c <= 9'b101110;
				8'b1000101: c <= 9'b100101000;
				8'b1011001: c <= 9'b11000;
				8'b110100: c <= 9'b10101001;
				8'b1111001: c <= 9'b111111010;
				8'b1110001: c <= 9'b101000101;
				8'b1001111: c <= 9'b100010100;
				8'b1100101: c <= 9'b101110101;
				8'b1111110: c <= 9'b10010001;
				8'b1111100: c <= 9'b1000010;
				8'b1010110: c <= 9'b110011011;
				8'b110010: c <= 9'b110100101;
				8'b1101101: c <= 9'b11001001;
				8'b100011: c <= 9'b1001;
				8'b1110101: c <= 9'b1000100;
				8'b1111101: c <= 9'b1010101;
				8'b101001: c <= 9'b111001110;
				8'b1010010: c <= 9'b101000011;
				8'b1011000: c <= 9'b111000010;
				8'b101110: c <= 9'b10100;
				8'b1000001: c <= 9'b100101110;
				default: c <= 9'b0;
			endcase
			9'b1111000 : case(di)
				8'b1000011: c <= 9'b110000110;
				8'b101000: c <= 9'b10001101;
				8'b111010: c <= 9'b11111100;
				8'b110110: c <= 9'b100011001;
				8'b1100100: c <= 9'b11001;
				8'b1000000: c <= 9'b110101011;
				8'b1110110: c <= 9'b1;
				8'b100101: c <= 9'b10111010;
				8'b101111: c <= 9'b100101000;
				8'b100110: c <= 9'b1111011;
				8'b1100011: c <= 9'b100000110;
				8'b1001000: c <= 9'b101010010;
				8'b111000: c <= 9'b111000101;
				8'b110001: c <= 9'b100000000;
				8'b1010111: c <= 9'b11010111;
				8'b1001110: c <= 9'b1100001;
				8'b1101010: c <= 9'b1000000;
				8'b1001001: c <= 9'b110001111;
				8'b1100000: c <= 9'b11101001;
				8'b110111: c <= 9'b111111110;
				8'b1011101: c <= 9'b100001101;
				8'b1011011: c <= 9'b101101000;
				8'b111001: c <= 9'b111001;
				8'b1001010: c <= 9'b100101101;
				8'b110011: c <= 9'b11100010;
				8'b1101100: c <= 9'b10100010;
				8'b1110111: c <= 9'b1100100;
				8'b101011: c <= 9'b11011000;
				8'b1101011: c <= 9'b10011010;
				8'b111100: c <= 9'b101000010;
				8'b1000111: c <= 9'b10110111;
				8'b1011111: c <= 9'b11100111;
				8'b1110100: c <= 9'b100110000;
				8'b101101: c <= 9'b101100001;
				8'b1010011: c <= 9'b10011000;
				8'b1100001: c <= 9'b10111101;
				8'b110101: c <= 9'b100111111;
				8'b1000100: c <= 9'b111101000;
				8'b1010001: c <= 9'b111110110;
				8'b1010100: c <= 9'b110100001;
				8'b1100110: c <= 9'b110010001;
				8'b101010: c <= 9'b100111101;
				8'b1011110: c <= 9'b111100;
				8'b1100111: c <= 9'b110110011;
				8'b1011010: c <= 9'b110001;
				8'b1000010: c <= 9'b100011100;
				8'b111101: c <= 9'b110010110;
				8'b110000: c <= 9'b100110111;
				8'b111110: c <= 9'b11100101;
				8'b1100010: c <= 9'b111001100;
				8'b1110000: c <= 9'b101101110;
				8'b1101001: c <= 9'b111011110;
				8'b1110011: c <= 9'b111011001;
				8'b1001100: c <= 9'b110101110;
				8'b100001: c <= 9'b1000001;
				8'b1000110: c <= 9'b111111110;
				8'b1110010: c <= 9'b111011010;
				8'b1010000: c <= 9'b10111110;
				8'b1111010: c <= 9'b100101100;
				8'b1010101: c <= 9'b100101011;
				8'b111011: c <= 9'b100011011;
				8'b1001101: c <= 9'b1100100;
				8'b111111: c <= 9'b111001;
				8'b1101110: c <= 9'b1000001;
				8'b1111011: c <= 9'b110011110;
				8'b1001011: c <= 9'b111011010;
				8'b1101111: c <= 9'b1111010;
				8'b1101000: c <= 9'b110101101;
				8'b101100: c <= 9'b111111001;
				8'b100100: c <= 9'b111000011;
				8'b1111000: c <= 9'b100100001;
				8'b1000101: c <= 9'b110011011;
				8'b1011001: c <= 9'b1000100;
				8'b110100: c <= 9'b110;
				8'b1111001: c <= 9'b111111101;
				8'b1110001: c <= 9'b1010111;
				8'b1001111: c <= 9'b100001110;
				8'b1100101: c <= 9'b100111110;
				8'b1111110: c <= 9'b11010000;
				8'b1111100: c <= 9'b11100001;
				8'b1010110: c <= 9'b1000100;
				8'b110010: c <= 9'b10011000;
				8'b1101101: c <= 9'b11110011;
				8'b100011: c <= 9'b11001111;
				8'b1110101: c <= 9'b110000;
				8'b1111101: c <= 9'b100100001;
				8'b101001: c <= 9'b1011111;
				8'b1010010: c <= 9'b111001111;
				8'b1011000: c <= 9'b10111110;
				8'b101110: c <= 9'b100000011;
				8'b1000001: c <= 9'b110000101;
				default: c <= 9'b0;
			endcase
			9'b10010101 : case(di)
				8'b1000011: c <= 9'b100011;
				8'b101000: c <= 9'b100011;
				8'b111010: c <= 9'b1100100;
				8'b110110: c <= 9'b110001;
				8'b1100100: c <= 9'b11100111;
				8'b1000000: c <= 9'b110101111;
				8'b1110110: c <= 9'b101100110;
				8'b100101: c <= 9'b110011011;
				8'b101111: c <= 9'b101010001;
				8'b100110: c <= 9'b100101111;
				8'b1100011: c <= 9'b110111001;
				8'b1001000: c <= 9'b110001010;
				8'b111000: c <= 9'b100010101;
				8'b110001: c <= 9'b110011111;
				8'b1010111: c <= 9'b101000100;
				8'b1001110: c <= 9'b100001;
				8'b1101010: c <= 9'b111010000;
				8'b1001001: c <= 9'b1111000;
				8'b1100000: c <= 9'b111101111;
				8'b110111: c <= 9'b101110001;
				8'b1011101: c <= 9'b10000111;
				8'b1011011: c <= 9'b11011001;
				8'b111001: c <= 9'b1100000;
				8'b1001010: c <= 9'b11111011;
				8'b110011: c <= 9'b101100010;
				8'b1101100: c <= 9'b110100111;
				8'b1110111: c <= 9'b10110111;
				8'b101011: c <= 9'b100111000;
				8'b1101011: c <= 9'b100010;
				8'b111100: c <= 9'b111100;
				8'b1000111: c <= 9'b110001001;
				8'b1011111: c <= 9'b11010111;
				8'b1110100: c <= 9'b100011001;
				8'b101101: c <= 9'b111110011;
				8'b1010011: c <= 9'b1000;
				8'b1100001: c <= 9'b100101;
				8'b110101: c <= 9'b11010011;
				8'b1000100: c <= 9'b101010;
				8'b1010001: c <= 9'b1101110;
				8'b1010100: c <= 9'b100101100;
				8'b1100110: c <= 9'b100111111;
				8'b101010: c <= 9'b101000100;
				8'b1011110: c <= 9'b110110101;
				8'b1100111: c <= 9'b10001110;
				8'b1011010: c <= 9'b100011011;
				8'b1000010: c <= 9'b110110000;
				8'b111101: c <= 9'b11001111;
				8'b110000: c <= 9'b10000110;
				8'b111110: c <= 9'b1000010;
				8'b1100010: c <= 9'b101111001;
				8'b1110000: c <= 9'b1101001;
				8'b1101001: c <= 9'b11110011;
				8'b1110011: c <= 9'b101011;
				8'b1001100: c <= 9'b110000111;
				8'b100001: c <= 9'b10011;
				8'b1000110: c <= 9'b1010110;
				8'b1110010: c <= 9'b1000;
				8'b1010000: c <= 9'b110000011;
				8'b1111010: c <= 9'b11011110;
				8'b1010101: c <= 9'b101110100;
				8'b111011: c <= 9'b100111111;
				8'b1001101: c <= 9'b100100011;
				8'b111111: c <= 9'b111011;
				8'b1101110: c <= 9'b101;
				8'b1111011: c <= 9'b1011111;
				8'b1001011: c <= 9'b1101110;
				8'b1101111: c <= 9'b10001001;
				8'b1101000: c <= 9'b110110101;
				8'b101100: c <= 9'b1010011;
				8'b100100: c <= 9'b111001000;
				8'b1111000: c <= 9'b101011110;
				8'b1000101: c <= 9'b1111010;
				8'b1011001: c <= 9'b100000001;
				8'b110100: c <= 9'b101001011;
				8'b1111001: c <= 9'b1110010;
				8'b1110001: c <= 9'b1011111;
				8'b1001111: c <= 9'b1110000;
				8'b1100101: c <= 9'b100011001;
				8'b1111110: c <= 9'b11101101;
				8'b1111100: c <= 9'b10101100;
				8'b1010110: c <= 9'b110000110;
				8'b110010: c <= 9'b101010011;
				8'b1101101: c <= 9'b101000011;
				8'b100011: c <= 9'b101101;
				8'b1110101: c <= 9'b11111011;
				8'b1111101: c <= 9'b1101010;
				8'b101001: c <= 9'b101000110;
				8'b1010010: c <= 9'b11001001;
				8'b1011000: c <= 9'b101110111;
				8'b101110: c <= 9'b111100100;
				8'b1000001: c <= 9'b10011101;
				default: c <= 9'b0;
			endcase
			9'b101110010 : case(di)
				8'b1000011: c <= 9'b10111;
				8'b101000: c <= 9'b10101000;
				8'b111010: c <= 9'b101111000;
				8'b110110: c <= 9'b11000010;
				8'b1100100: c <= 9'b100100111;
				8'b1000000: c <= 9'b111001101;
				8'b1110110: c <= 9'b10110101;
				8'b100101: c <= 9'b101000010;
				8'b101111: c <= 9'b111100011;
				8'b100110: c <= 9'b111010001;
				8'b1100011: c <= 9'b10010011;
				8'b1001000: c <= 9'b110010010;
				8'b111000: c <= 9'b110101001;
				8'b110001: c <= 9'b10011111;
				8'b1010111: c <= 9'b110001101;
				8'b1001110: c <= 9'b110010001;
				8'b1101010: c <= 9'b100000001;
				8'b1001001: c <= 9'b110011001;
				8'b1100000: c <= 9'b1110011;
				8'b110111: c <= 9'b10000;
				8'b1011101: c <= 9'b100001100;
				8'b1011011: c <= 9'b101100110;
				8'b111001: c <= 9'b101110010;
				8'b1001010: c <= 9'b1110011;
				8'b110011: c <= 9'b110000;
				8'b1101100: c <= 9'b11000;
				8'b1110111: c <= 9'b11001100;
				8'b101011: c <= 9'b11011100;
				8'b1101011: c <= 9'b100011000;
				8'b111100: c <= 9'b111000101;
				8'b1000111: c <= 9'b110001010;
				8'b1011111: c <= 9'b100110011;
				8'b1110100: c <= 9'b111111000;
				8'b101101: c <= 9'b101001;
				8'b1010011: c <= 9'b111001;
				8'b1100001: c <= 9'b10001110;
				8'b110101: c <= 9'b110010;
				8'b1000100: c <= 9'b10000111;
				8'b1010001: c <= 9'b10011100;
				8'b1010100: c <= 9'b101100100;
				8'b1100110: c <= 9'b110000101;
				8'b101010: c <= 9'b101001111;
				8'b1011110: c <= 9'b1100101;
				8'b1100111: c <= 9'b111110000;
				8'b1011010: c <= 9'b10101101;
				8'b1000010: c <= 9'b110111100;
				8'b111101: c <= 9'b10001110;
				8'b110000: c <= 9'b1100011;
				8'b111110: c <= 9'b101111000;
				8'b1100010: c <= 9'b1011010;
				8'b1110000: c <= 9'b110100000;
				8'b1101001: c <= 9'b1100111;
				8'b1110011: c <= 9'b111100101;
				8'b1001100: c <= 9'b110101001;
				8'b100001: c <= 9'b110000111;
				8'b1000110: c <= 9'b11110;
				8'b1110010: c <= 9'b110011011;
				8'b1010000: c <= 9'b11110100;
				8'b1111010: c <= 9'b110101111;
				8'b1010101: c <= 9'b101100100;
				8'b111011: c <= 9'b10000111;
				8'b1001101: c <= 9'b1111101;
				8'b111111: c <= 9'b100000001;
				8'b1101110: c <= 9'b10011111;
				8'b1111011: c <= 9'b111011001;
				8'b1001011: c <= 9'b11001100;
				8'b1101111: c <= 9'b100010101;
				8'b1101000: c <= 9'b110111011;
				8'b101100: c <= 9'b10101;
				8'b100100: c <= 9'b110101011;
				8'b1111000: c <= 9'b1001010;
				8'b1000101: c <= 9'b1010010;
				8'b1011001: c <= 9'b101100010;
				8'b110100: c <= 9'b11100011;
				8'b1111001: c <= 9'b10010011;
				8'b1110001: c <= 9'b1100101;
				8'b1001111: c <= 9'b111001;
				8'b1100101: c <= 9'b101110011;
				8'b1111110: c <= 9'b110100111;
				8'b1111100: c <= 9'b111001;
				8'b1010110: c <= 9'b10001101;
				8'b110010: c <= 9'b1000010;
				8'b1101101: c <= 9'b111101001;
				8'b100011: c <= 9'b10010110;
				8'b1110101: c <= 9'b101011001;
				8'b1111101: c <= 9'b101011001;
				8'b101001: c <= 9'b111110001;
				8'b1010010: c <= 9'b110100000;
				8'b1011000: c <= 9'b10000;
				8'b101110: c <= 9'b11101;
				8'b1000001: c <= 9'b11000010;
				default: c <= 9'b0;
			endcase
			9'b11100010 : case(di)
				8'b1000011: c <= 9'b100000101;
				8'b101000: c <= 9'b101101101;
				8'b111010: c <= 9'b11000010;
				8'b110110: c <= 9'b111000100;
				8'b1100100: c <= 9'b110000110;
				8'b1000000: c <= 9'b101110;
				8'b1110110: c <= 9'b100010100;
				8'b100101: c <= 9'b110001;
				8'b101111: c <= 9'b111000101;
				8'b100110: c <= 9'b110001001;
				8'b1100011: c <= 9'b100000100;
				8'b1001000: c <= 9'b11011110;
				8'b111000: c <= 9'b1111010;
				8'b110001: c <= 9'b11010001;
				8'b1010111: c <= 9'b11010101;
				8'b1001110: c <= 9'b11001011;
				8'b1101010: c <= 9'b11100111;
				8'b1001001: c <= 9'b11010111;
				8'b1100000: c <= 9'b11100101;
				8'b110111: c <= 9'b1111000;
				8'b1011101: c <= 9'b101010110;
				8'b1011011: c <= 9'b101100;
				8'b111001: c <= 9'b110010;
				8'b1001010: c <= 9'b101100011;
				8'b110011: c <= 9'b101010110;
				8'b1101100: c <= 9'b100110100;
				8'b1110111: c <= 9'b10111111;
				8'b101011: c <= 9'b111111001;
				8'b1101011: c <= 9'b100100011;
				8'b111100: c <= 9'b10110001;
				8'b1000111: c <= 9'b1000001;
				8'b1011111: c <= 9'b1000;
				8'b1110100: c <= 9'b10011101;
				8'b101101: c <= 9'b11110;
				8'b1010011: c <= 9'b11011110;
				8'b1100001: c <= 9'b100110101;
				8'b110101: c <= 9'b11110110;
				8'b1000100: c <= 9'b111100000;
				8'b1010001: c <= 9'b101110110;
				8'b1010100: c <= 9'b10110011;
				8'b1100110: c <= 9'b110100000;
				8'b101010: c <= 9'b1001111;
				8'b1011110: c <= 9'b100111001;
				8'b1100111: c <= 9'b1101110;
				8'b1011010: c <= 9'b101100111;
				8'b1000010: c <= 9'b1110111;
				8'b111101: c <= 9'b100011000;
				8'b110000: c <= 9'b1100001;
				8'b111110: c <= 9'b110101010;
				8'b1100010: c <= 9'b11100110;
				8'b1110000: c <= 9'b11111100;
				8'b1101001: c <= 9'b10101110;
				8'b1110011: c <= 9'b111010010;
				8'b1001100: c <= 9'b111000101;
				8'b100001: c <= 9'b11010011;
				8'b1000110: c <= 9'b11100001;
				8'b1110010: c <= 9'b111100110;
				8'b1010000: c <= 9'b110001;
				8'b1111010: c <= 9'b111101101;
				8'b1010101: c <= 9'b10000111;
				8'b111011: c <= 9'b111101101;
				8'b1001101: c <= 9'b110110;
				8'b111111: c <= 9'b100111001;
				8'b1101110: c <= 9'b101111001;
				8'b1111011: c <= 9'b110001001;
				8'b1001011: c <= 9'b111011;
				8'b1101111: c <= 9'b10100100;
				8'b1101000: c <= 9'b11100101;
				8'b101100: c <= 9'b11001011;
				8'b100100: c <= 9'b10000110;
				8'b1111000: c <= 9'b11111;
				8'b1000101: c <= 9'b1010111;
				8'b1011001: c <= 9'b111100101;
				8'b110100: c <= 9'b10011100;
				8'b1111001: c <= 9'b1111101;
				8'b1110001: c <= 9'b110011;
				8'b1001111: c <= 9'b11;
				8'b1100101: c <= 9'b101001010;
				8'b1111110: c <= 9'b100011111;
				8'b1111100: c <= 9'b100000010;
				8'b1010110: c <= 9'b101101101;
				8'b110010: c <= 9'b100011011;
				8'b1101101: c <= 9'b100101111;
				8'b100011: c <= 9'b101101;
				8'b1110101: c <= 9'b11101011;
				8'b1111101: c <= 9'b110010;
				8'b101001: c <= 9'b101100010;
				8'b1010010: c <= 9'b110011;
				8'b1011000: c <= 9'b100011011;
				8'b101110: c <= 9'b111001010;
				8'b1000001: c <= 9'b110000111;
				default: c <= 9'b0;
			endcase
			9'b110111000 : case(di)
				8'b1000011: c <= 9'b11001100;
				8'b101000: c <= 9'b10011101;
				8'b111010: c <= 9'b111010;
				8'b110110: c <= 9'b11011010;
				8'b1100100: c <= 9'b111001000;
				8'b1000000: c <= 9'b10011000;
				8'b1110110: c <= 9'b110000101;
				8'b100101: c <= 9'b10101100;
				8'b101111: c <= 9'b100101;
				8'b100110: c <= 9'b111011110;
				8'b1100011: c <= 9'b110111000;
				8'b1001000: c <= 9'b110001101;
				8'b111000: c <= 9'b111111010;
				8'b110001: c <= 9'b111100100;
				8'b1010111: c <= 9'b11000110;
				8'b1001110: c <= 9'b1001100;
				8'b1101010: c <= 9'b110101111;
				8'b1001001: c <= 9'b111100;
				8'b1100000: c <= 9'b101010001;
				8'b110111: c <= 9'b111010;
				8'b1011101: c <= 9'b10001000;
				8'b1011011: c <= 9'b100100110;
				8'b111001: c <= 9'b111011111;
				8'b1001010: c <= 9'b1011011;
				8'b110011: c <= 9'b100010010;
				8'b1101100: c <= 9'b10000001;
				8'b1110111: c <= 9'b111101100;
				8'b101011: c <= 9'b10100000;
				8'b1101011: c <= 9'b10101;
				8'b111100: c <= 9'b10011101;
				8'b1000111: c <= 9'b1101000;
				8'b1011111: c <= 9'b110101010;
				8'b1110100: c <= 9'b101001;
				8'b101101: c <= 9'b101001000;
				8'b1010011: c <= 9'b11;
				8'b1100001: c <= 9'b1100101;
				8'b110101: c <= 9'b1001001;
				8'b1000100: c <= 9'b10110011;
				8'b1010001: c <= 9'b11011001;
				8'b1010100: c <= 9'b110100110;
				8'b1100110: c <= 9'b1011011;
				8'b101010: c <= 9'b1100010;
				8'b1011110: c <= 9'b11110101;
				8'b1100111: c <= 9'b100001010;
				8'b1011010: c <= 9'b1111101;
				8'b1000010: c <= 9'b10010001;
				8'b111101: c <= 9'b101110001;
				8'b110000: c <= 9'b1110000;
				8'b111110: c <= 9'b10000;
				8'b1100010: c <= 9'b10011010;
				8'b1110000: c <= 9'b1001000;
				8'b1101001: c <= 9'b100110110;
				8'b1110011: c <= 9'b1000001;
				8'b1001100: c <= 9'b1110;
				8'b100001: c <= 9'b100010100;
				8'b1000110: c <= 9'b11111001;
				8'b1110010: c <= 9'b111000100;
				8'b1010000: c <= 9'b10000101;
				8'b1111010: c <= 9'b101111010;
				8'b1010101: c <= 9'b111001111;
				8'b111011: c <= 9'b11000001;
				8'b1001101: c <= 9'b10101000;
				8'b111111: c <= 9'b11111010;
				8'b1101110: c <= 9'b1010110;
				8'b1111011: c <= 9'b1010011;
				8'b1001011: c <= 9'b1010000;
				8'b1101111: c <= 9'b111011;
				8'b1101000: c <= 9'b11101011;
				8'b101100: c <= 9'b11101101;
				8'b100100: c <= 9'b11000100;
				8'b1111000: c <= 9'b1111000;
				8'b1000101: c <= 9'b110100011;
				8'b1011001: c <= 9'b110011001;
				8'b110100: c <= 9'b110101001;
				8'b1111001: c <= 9'b111000100;
				8'b1110001: c <= 9'b101101100;
				8'b1001111: c <= 9'b111110110;
				8'b1100101: c <= 9'b100010101;
				8'b1111110: c <= 9'b110;
				8'b1111100: c <= 9'b111110110;
				8'b1010110: c <= 9'b10010100;
				8'b110010: c <= 9'b100100010;
				8'b1101101: c <= 9'b11110101;
				8'b100011: c <= 9'b110111110;
				8'b1110101: c <= 9'b1111111;
				8'b1111101: c <= 9'b111000;
				8'b101001: c <= 9'b1101010;
				8'b1010010: c <= 9'b10001101;
				8'b1011000: c <= 9'b110100111;
				8'b101110: c <= 9'b1100000;
				8'b1000001: c <= 9'b111110101;
				default: c <= 9'b0;
			endcase
			9'b111111000 : case(di)
				8'b1000011: c <= 9'b11010100;
				8'b101000: c <= 9'b10010100;
				8'b111010: c <= 9'b111100110;
				8'b110110: c <= 9'b1111000;
				8'b1100100: c <= 9'b100110100;
				8'b1000000: c <= 9'b1001010;
				8'b1110110: c <= 9'b11111101;
				8'b100101: c <= 9'b1001011;
				8'b101111: c <= 9'b1100001;
				8'b100110: c <= 9'b11011011;
				8'b1100011: c <= 9'b100101010;
				8'b1001000: c <= 9'b111001110;
				8'b111000: c <= 9'b110011101;
				8'b110001: c <= 9'b101011011;
				8'b1010111: c <= 9'b1110;
				8'b1001110: c <= 9'b110001101;
				8'b1101010: c <= 9'b11011100;
				8'b1001001: c <= 9'b100001010;
				8'b1100000: c <= 9'b11001110;
				8'b110111: c <= 9'b10000111;
				8'b1011101: c <= 9'b110101111;
				8'b1011011: c <= 9'b100001110;
				8'b111001: c <= 9'b10001000;
				8'b1001010: c <= 9'b110110110;
				8'b110011: c <= 9'b1011011;
				8'b1101100: c <= 9'b11110111;
				8'b1110111: c <= 9'b1010001;
				8'b101011: c <= 9'b111101000;
				8'b1101011: c <= 9'b110011110;
				8'b111100: c <= 9'b10101001;
				8'b1000111: c <= 9'b10101000;
				8'b1011111: c <= 9'b1111111;
				8'b1110100: c <= 9'b10011101;
				8'b101101: c <= 9'b111111011;
				8'b1010011: c <= 9'b101011;
				8'b1100001: c <= 9'b10011000;
				8'b110101: c <= 9'b111001100;
				8'b1000100: c <= 9'b110011101;
				8'b1010001: c <= 9'b1111100;
				8'b1010100: c <= 9'b100100011;
				8'b1100110: c <= 9'b10001011;
				8'b101010: c <= 9'b100111110;
				8'b1011110: c <= 9'b11100100;
				8'b1100111: c <= 9'b1101110;
				8'b1011010: c <= 9'b11100001;
				8'b1000010: c <= 9'b1011001;
				8'b111101: c <= 9'b111010000;
				8'b110000: c <= 9'b101110100;
				8'b111110: c <= 9'b110100110;
				8'b1100010: c <= 9'b1000010;
				8'b1110000: c <= 9'b110101001;
				8'b1101001: c <= 9'b111001101;
				8'b1110011: c <= 9'b111100100;
				8'b1001100: c <= 9'b11101011;
				8'b100001: c <= 9'b101100110;
				8'b1000110: c <= 9'b110011000;
				8'b1110010: c <= 9'b100010100;
				8'b1010000: c <= 9'b101010;
				8'b1111010: c <= 9'b100111;
				8'b1010101: c <= 9'b101;
				8'b111011: c <= 9'b101101010;
				8'b1001101: c <= 9'b10010111;
				8'b111111: c <= 9'b110011000;
				8'b1101110: c <= 9'b1001110;
				8'b1111011: c <= 9'b110011110;
				8'b1001011: c <= 9'b100110101;
				8'b1101111: c <= 9'b101001100;
				8'b1101000: c <= 9'b100100;
				8'b101100: c <= 9'b110100000;
				8'b100100: c <= 9'b1011100;
				8'b1111000: c <= 9'b101011110;
				8'b1000101: c <= 9'b10101;
				8'b1011001: c <= 9'b11000;
				8'b110100: c <= 9'b10010;
				8'b1111001: c <= 9'b10100010;
				8'b1110001: c <= 9'b110000101;
				8'b1001111: c <= 9'b10111011;
				8'b1100101: c <= 9'b11101011;
				8'b1111110: c <= 9'b101010011;
				8'b1111100: c <= 9'b10000000;
				8'b1010110: c <= 9'b11111001;
				8'b110010: c <= 9'b100100111;
				8'b1101101: c <= 9'b101010001;
				8'b100011: c <= 9'b1101100;
				8'b1110101: c <= 9'b10011;
				8'b1111101: c <= 9'b110100000;
				8'b101001: c <= 9'b110100;
				8'b1010010: c <= 9'b10;
				8'b1011000: c <= 9'b110100101;
				8'b101110: c <= 9'b111010110;
				8'b1000001: c <= 9'b111100100;
				default: c <= 9'b0;
			endcase
			9'b100101 : case(di)
				8'b1000011: c <= 9'b1111010;
				8'b101000: c <= 9'b101000;
				8'b111010: c <= 9'b110100011;
				8'b110110: c <= 9'b111101010;
				8'b1100100: c <= 9'b100011010;
				8'b1000000: c <= 9'b111010;
				8'b1110110: c <= 9'b100000101;
				8'b100101: c <= 9'b10010101;
				8'b101111: c <= 9'b111111000;
				8'b100110: c <= 9'b110100001;
				8'b1100011: c <= 9'b110101101;
				8'b1001000: c <= 9'b11001101;
				8'b111000: c <= 9'b110001100;
				8'b110001: c <= 9'b101111000;
				8'b1010111: c <= 9'b1101111;
				8'b1001110: c <= 9'b100001101;
				8'b1101010: c <= 9'b1011111;
				8'b1001001: c <= 9'b101101100;
				8'b1100000: c <= 9'b101100001;
				8'b110111: c <= 9'b100111001;
				8'b1011101: c <= 9'b101101111;
				8'b1011011: c <= 9'b100110111;
				8'b111001: c <= 9'b100010;
				8'b1001010: c <= 9'b11100100;
				8'b110011: c <= 9'b101001111;
				8'b1101100: c <= 9'b100001;
				8'b1110111: c <= 9'b111001000;
				8'b101011: c <= 9'b110010011;
				8'b1101011: c <= 9'b10111;
				8'b111100: c <= 9'b11111010;
				8'b1000111: c <= 9'b101110110;
				8'b1011111: c <= 9'b111001;
				8'b1110100: c <= 9'b1110100;
				8'b101101: c <= 9'b11011101;
				8'b1010011: c <= 9'b100000000;
				8'b1100001: c <= 9'b10100;
				8'b110101: c <= 9'b101100001;
				8'b1000100: c <= 9'b110011011;
				8'b1010001: c <= 9'b1110001;
				8'b1010100: c <= 9'b100000100;
				8'b1100110: c <= 9'b1111000;
				8'b101010: c <= 9'b100100;
				8'b1011110: c <= 9'b11011011;
				8'b1100111: c <= 9'b100110000;
				8'b1011010: c <= 9'b1010011;
				8'b1000010: c <= 9'b101000110;
				8'b111101: c <= 9'b11011010;
				8'b110000: c <= 9'b110001100;
				8'b111110: c <= 9'b111111001;
				8'b1100010: c <= 9'b101110000;
				8'b1110000: c <= 9'b111011;
				8'b1101001: c <= 9'b1101010;
				8'b1110011: c <= 9'b110011;
				8'b1001100: c <= 9'b100110011;
				8'b100001: c <= 9'b110000101;
				8'b1000110: c <= 9'b111000011;
				8'b1110010: c <= 9'b101010011;
				8'b1010000: c <= 9'b110101100;
				8'b1111010: c <= 9'b111001010;
				8'b1010101: c <= 9'b111001010;
				8'b111011: c <= 9'b11111000;
				8'b1001101: c <= 9'b100001100;
				8'b111111: c <= 9'b1101101;
				8'b1101110: c <= 9'b1001001;
				8'b1111011: c <= 9'b11001001;
				8'b1001011: c <= 9'b10011;
				8'b1101111: c <= 9'b1101111;
				8'b1101000: c <= 9'b1100001;
				8'b101100: c <= 9'b10000011;
				8'b100100: c <= 9'b110010111;
				8'b1111000: c <= 9'b10001101;
				8'b1000101: c <= 9'b100101110;
				8'b1011001: c <= 9'b10001100;
				8'b110100: c <= 9'b111001010;
				8'b1111001: c <= 9'b1101001;
				8'b1110001: c <= 9'b1101111;
				8'b1001111: c <= 9'b1000111;
				8'b1100101: c <= 9'b111111101;
				8'b1111110: c <= 9'b11111011;
				8'b1111100: c <= 9'b10010001;
				8'b1010110: c <= 9'b110110101;
				8'b110010: c <= 9'b111111010;
				8'b1101101: c <= 9'b101101101;
				8'b100011: c <= 9'b111000;
				8'b1110101: c <= 9'b11011000;
				8'b1111101: c <= 9'b101011011;
				8'b101001: c <= 9'b10011010;
				8'b1010010: c <= 9'b100100111;
				8'b1011000: c <= 9'b111110110;
				8'b101110: c <= 9'b10001111;
				8'b1000001: c <= 9'b100110110;
				default: c <= 9'b0;
			endcase
			9'b100000100 : case(di)
				8'b1000011: c <= 9'b10111010;
				8'b101000: c <= 9'b10110010;
				8'b111010: c <= 9'b110101;
				8'b110110: c <= 9'b11011010;
				8'b1100100: c <= 9'b101001011;
				8'b1000000: c <= 9'b11101100;
				8'b1110110: c <= 9'b10111010;
				8'b100101: c <= 9'b1001000;
				8'b101111: c <= 9'b1001000;
				8'b100110: c <= 9'b1110111;
				8'b1100011: c <= 9'b101001100;
				8'b1001000: c <= 9'b110100100;
				8'b111000: c <= 9'b1000011;
				8'b110001: c <= 9'b11001100;
				8'b1010111: c <= 9'b10101001;
				8'b1001110: c <= 9'b10001011;
				8'b1101010: c <= 9'b1001010;
				8'b1001001: c <= 9'b100100010;
				8'b1100000: c <= 9'b111001010;
				8'b110111: c <= 9'b111010100;
				8'b1011101: c <= 9'b101000111;
				8'b1011011: c <= 9'b111;
				8'b111001: c <= 9'b1001;
				8'b1001010: c <= 9'b111000010;
				8'b110011: c <= 9'b101101011;
				8'b1101100: c <= 9'b100011100;
				8'b1110111: c <= 9'b111001;
				8'b101011: c <= 9'b101010110;
				8'b1101011: c <= 9'b100010010;
				8'b111100: c <= 9'b100100101;
				8'b1000111: c <= 9'b1100111;
				8'b1011111: c <= 9'b101110101;
				8'b1110100: c <= 9'b11101000;
				8'b101101: c <= 9'b100000101;
				8'b1010011: c <= 9'b101001;
				8'b1100001: c <= 9'b100001;
				8'b110101: c <= 9'b10001111;
				8'b1000100: c <= 9'b101101110;
				8'b1010001: c <= 9'b110110111;
				8'b1010100: c <= 9'b11111001;
				8'b1100110: c <= 9'b110100110;
				8'b101010: c <= 9'b1110101;
				8'b1011110: c <= 9'b1001111;
				8'b1100111: c <= 9'b101001100;
				8'b1011010: c <= 9'b110111010;
				8'b1000010: c <= 9'b10000011;
				8'b111101: c <= 9'b110000;
				8'b110000: c <= 9'b11110101;
				8'b111110: c <= 9'b11101101;
				8'b1100010: c <= 9'b11111010;
				8'b1110000: c <= 9'b110001;
				8'b1101001: c <= 9'b10110101;
				8'b1110011: c <= 9'b11100001;
				8'b1001100: c <= 9'b100101010;
				8'b100001: c <= 9'b110001101;
				8'b1000110: c <= 9'b11011;
				8'b1110010: c <= 9'b1000;
				8'b1010000: c <= 9'b111001000;
				8'b1111010: c <= 9'b110010010;
				8'b1010101: c <= 9'b110010010;
				8'b111011: c <= 9'b101111010;
				8'b1001101: c <= 9'b10010100;
				8'b111111: c <= 9'b110010001;
				8'b1101110: c <= 9'b10100000;
				8'b1111011: c <= 9'b1000;
				8'b1001011: c <= 9'b10010101;
				8'b1101111: c <= 9'b110001101;
				8'b1101000: c <= 9'b110011001;
				8'b101100: c <= 9'b111010;
				8'b100100: c <= 9'b10111110;
				8'b1111000: c <= 9'b111001000;
				8'b1000101: c <= 9'b10011011;
				8'b1011001: c <= 9'b110111010;
				8'b110100: c <= 9'b1111100;
				8'b1111001: c <= 9'b10100110;
				8'b1110001: c <= 9'b10111010;
				8'b1001111: c <= 9'b11011101;
				8'b1100101: c <= 9'b11110001;
				8'b1111110: c <= 9'b1000100;
				8'b1111100: c <= 9'b1100;
				8'b1010110: c <= 9'b101000;
				8'b110010: c <= 9'b1000011;
				8'b1101101: c <= 9'b10010110;
				8'b100011: c <= 9'b101100100;
				8'b1110101: c <= 9'b100111;
				8'b1111101: c <= 9'b11111011;
				8'b101001: c <= 9'b100101111;
				8'b1010010: c <= 9'b111110011;
				8'b1011000: c <= 9'b11100;
				8'b101110: c <= 9'b101110000;
				8'b1000001: c <= 9'b111111110;
				default: c <= 9'b0;
			endcase
			9'b11100 : case(di)
				8'b1000011: c <= 9'b10010100;
				8'b101000: c <= 9'b101101100;
				8'b111010: c <= 9'b10110010;
				8'b110110: c <= 9'b11111100;
				8'b1100100: c <= 9'b111101001;
				8'b1000000: c <= 9'b101101001;
				8'b1110110: c <= 9'b110110010;
				8'b100101: c <= 9'b110110101;
				8'b101111: c <= 9'b101111001;
				8'b100110: c <= 9'b1000111;
				8'b1100011: c <= 9'b110110010;
				8'b1001000: c <= 9'b101000001;
				8'b111000: c <= 9'b101101100;
				8'b110001: c <= 9'b101110111;
				8'b1010111: c <= 9'b111010010;
				8'b1001110: c <= 9'b111111;
				8'b1101010: c <= 9'b10011101;
				8'b1001001: c <= 9'b11100001;
				8'b1100000: c <= 9'b101000011;
				8'b110111: c <= 9'b11001101;
				8'b1011101: c <= 9'b100011101;
				8'b1011011: c <= 9'b111010;
				8'b111001: c <= 9'b110111001;
				8'b1001010: c <= 9'b10010101;
				8'b110011: c <= 9'b100110110;
				8'b1101100: c <= 9'b11110101;
				8'b1110111: c <= 9'b110001001;
				8'b101011: c <= 9'b11110110;
				8'b1101011: c <= 9'b10001111;
				8'b111100: c <= 9'b11100010;
				8'b1000111: c <= 9'b11000010;
				8'b1011111: c <= 9'b110110010;
				8'b1110100: c <= 9'b101100111;
				8'b101101: c <= 9'b10010100;
				8'b1010011: c <= 9'b111110101;
				8'b1100001: c <= 9'b1000011;
				8'b110101: c <= 9'b11101;
				8'b1000100: c <= 9'b11101000;
				8'b1010001: c <= 9'b100010010;
				8'b1010100: c <= 9'b111111001;
				8'b1100110: c <= 9'b11010011;
				8'b101010: c <= 9'b11101;
				8'b1011110: c <= 9'b10011111;
				8'b1100111: c <= 9'b10001001;
				8'b1011010: c <= 9'b10000110;
				8'b1000010: c <= 9'b101101000;
				8'b111101: c <= 9'b1001101;
				8'b110000: c <= 9'b101011011;
				8'b111110: c <= 9'b111001110;
				8'b1100010: c <= 9'b10000000;
				8'b1110000: c <= 9'b111101100;
				8'b1101001: c <= 9'b110110000;
				8'b1110011: c <= 9'b110010111;
				8'b1001100: c <= 9'b1100000;
				8'b100001: c <= 9'b101011111;
				8'b1000110: c <= 9'b10000110;
				8'b1110010: c <= 9'b111110110;
				8'b1010000: c <= 9'b1111100;
				8'b1111010: c <= 9'b111111111;
				8'b1010101: c <= 9'b101011111;
				8'b111011: c <= 9'b110111000;
				8'b1001101: c <= 9'b1101111;
				8'b111111: c <= 9'b1000011;
				8'b1101110: c <= 9'b100100101;
				8'b1111011: c <= 9'b110011010;
				8'b1001011: c <= 9'b10101;
				8'b1101111: c <= 9'b1001110;
				8'b1101000: c <= 9'b1010000;
				8'b101100: c <= 9'b11001011;
				8'b100100: c <= 9'b11000100;
				8'b1111000: c <= 9'b111110000;
				8'b1000101: c <= 9'b100010110;
				8'b1011001: c <= 9'b11011;
				8'b110100: c <= 9'b100101;
				8'b1111001: c <= 9'b100100;
				8'b1110001: c <= 9'b11100100;
				8'b1001111: c <= 9'b110100;
				8'b1100101: c <= 9'b110101100;
				8'b1111110: c <= 9'b1100101;
				8'b1111100: c <= 9'b110110100;
				8'b1010110: c <= 9'b110000001;
				8'b110010: c <= 9'b11001;
				8'b1101101: c <= 9'b101011011;
				8'b100011: c <= 9'b111111001;
				8'b1110101: c <= 9'b10110100;
				8'b1111101: c <= 9'b111011110;
				8'b101001: c <= 9'b110011001;
				8'b1010010: c <= 9'b1100010;
				8'b1011000: c <= 9'b11111011;
				8'b101110: c <= 9'b101100011;
				8'b1000001: c <= 9'b110010110;
				default: c <= 9'b0;
			endcase
			9'b111000 : case(di)
				8'b1000011: c <= 9'b1001;
				8'b101000: c <= 9'b111011;
				8'b111010: c <= 9'b1001000;
				8'b110110: c <= 9'b100010011;
				8'b1100100: c <= 9'b101010100;
				8'b1000000: c <= 9'b1001101;
				8'b1110110: c <= 9'b100111101;
				8'b100101: c <= 9'b1110101;
				8'b101111: c <= 9'b1110011;
				8'b100110: c <= 9'b100011101;
				8'b1100011: c <= 9'b110001001;
				8'b1001000: c <= 9'b111111001;
				8'b111000: c <= 9'b101110110;
				8'b110001: c <= 9'b1001000;
				8'b1010111: c <= 9'b111100100;
				8'b1001110: c <= 9'b110010001;
				8'b1101010: c <= 9'b111001101;
				8'b1001001: c <= 9'b111110110;
				8'b1100000: c <= 9'b1101111;
				8'b110111: c <= 9'b10011;
				8'b1011101: c <= 9'b10110011;
				8'b1011011: c <= 9'b111110110;
				8'b111001: c <= 9'b100111100;
				8'b1001010: c <= 9'b101101001;
				8'b110011: c <= 9'b111101001;
				8'b1101100: c <= 9'b11011010;
				8'b1110111: c <= 9'b100100111;
				8'b101011: c <= 9'b101101011;
				8'b1101011: c <= 9'b111001001;
				8'b111100: c <= 9'b1010010;
				8'b1000111: c <= 9'b111001001;
				8'b1011111: c <= 9'b111000100;
				8'b1110100: c <= 9'b1010001;
				8'b101101: c <= 9'b111001001;
				8'b1010011: c <= 9'b11011100;
				8'b1100001: c <= 9'b11010100;
				8'b110101: c <= 9'b101100010;
				8'b1000100: c <= 9'b110000;
				8'b1010001: c <= 9'b1110010;
				8'b1010100: c <= 9'b1110;
				8'b1100110: c <= 9'b11001111;
				8'b101010: c <= 9'b110111110;
				8'b1011110: c <= 9'b110110000;
				8'b1100111: c <= 9'b10000001;
				8'b1011010: c <= 9'b111010100;
				8'b1000010: c <= 9'b100010000;
				8'b111101: c <= 9'b101101;
				8'b110000: c <= 9'b1010110;
				8'b111110: c <= 9'b101111110;
				8'b1100010: c <= 9'b10000000;
				8'b1110000: c <= 9'b111111111;
				8'b1101001: c <= 9'b110110101;
				8'b1110011: c <= 9'b11110001;
				8'b1001100: c <= 9'b110001001;
				8'b100001: c <= 9'b1101;
				8'b1000110: c <= 9'b10101110;
				8'b1110010: c <= 9'b11011101;
				8'b1010000: c <= 9'b1010111;
				8'b1111010: c <= 9'b11101011;
				8'b1010101: c <= 9'b10111110;
				8'b111011: c <= 9'b11010001;
				8'b1001101: c <= 9'b11010111;
				8'b111111: c <= 9'b101011;
				8'b1101110: c <= 9'b11110000;
				8'b1111011: c <= 9'b11100010;
				8'b1001011: c <= 9'b1001101;
				8'b1101111: c <= 9'b10111101;
				8'b1101000: c <= 9'b110011;
				8'b101100: c <= 9'b10000;
				8'b100100: c <= 9'b100111111;
				8'b1111000: c <= 9'b1101000;
				8'b1000101: c <= 9'b10100011;
				8'b1011001: c <= 9'b10000001;
				8'b110100: c <= 9'b110001100;
				8'b1111001: c <= 9'b101001111;
				8'b1110001: c <= 9'b110111;
				8'b1001111: c <= 9'b110001;
				8'b1100101: c <= 9'b10000110;
				8'b1111110: c <= 9'b11001;
				8'b1111100: c <= 9'b101010110;
				8'b1010110: c <= 9'b100010011;
				8'b110010: c <= 9'b1111010;
				8'b1101101: c <= 9'b11011001;
				8'b100011: c <= 9'b10000000;
				8'b1110101: c <= 9'b110101010;
				8'b1111101: c <= 9'b1011110;
				8'b101001: c <= 9'b10110100;
				8'b1010010: c <= 9'b110100000;
				8'b1011000: c <= 9'b1110;
				8'b101110: c <= 9'b101001;
				8'b1000001: c <= 9'b11011100;
				default: c <= 9'b0;
			endcase
			9'b100101000 : case(di)
				8'b1000011: c <= 9'b101101101;
				8'b101000: c <= 9'b111110001;
				8'b111010: c <= 9'b11100011;
				8'b110110: c <= 9'b111000101;
				8'b1100100: c <= 9'b11111;
				8'b1000000: c <= 9'b11011101;
				8'b1110110: c <= 9'b1111010;
				8'b100101: c <= 9'b110011;
				8'b101111: c <= 9'b11110101;
				8'b100110: c <= 9'b11111001;
				8'b1100011: c <= 9'b10111101;
				8'b1001000: c <= 9'b11100010;
				8'b111000: c <= 9'b111101;
				8'b110001: c <= 9'b1011;
				8'b1010111: c <= 9'b11110000;
				8'b1001110: c <= 9'b100100111;
				8'b1101010: c <= 9'b10010110;
				8'b1001001: c <= 9'b111111110;
				8'b1100000: c <= 9'b110;
				8'b110111: c <= 9'b111101110;
				8'b1011101: c <= 9'b11000001;
				8'b1011011: c <= 9'b100100111;
				8'b111001: c <= 9'b1101001;
				8'b1001010: c <= 9'b100101101;
				8'b110011: c <= 9'b101010111;
				8'b1101100: c <= 9'b100111001;
				8'b1110111: c <= 9'b1000011;
				8'b101011: c <= 9'b111100111;
				8'b1101011: c <= 9'b100010000;
				8'b111100: c <= 9'b11110110;
				8'b1000111: c <= 9'b111001010;
				8'b1011111: c <= 9'b110001111;
				8'b1110100: c <= 9'b10111110;
				8'b101101: c <= 9'b111011;
				8'b1010011: c <= 9'b101100010;
				8'b1100001: c <= 9'b101010101;
				8'b110101: c <= 9'b100010111;
				8'b1000100: c <= 9'b11101011;
				8'b1010001: c <= 9'b110011101;
				8'b1010100: c <= 9'b101011010;
				8'b1100110: c <= 9'b111000101;
				8'b101010: c <= 9'b11100000;
				8'b1011110: c <= 9'b10100100;
				8'b1100111: c <= 9'b111000111;
				8'b1011010: c <= 9'b11101100;
				8'b1000010: c <= 9'b10001010;
				8'b111101: c <= 9'b11000000;
				8'b110000: c <= 9'b10101101;
				8'b111110: c <= 9'b100001001;
				8'b1100010: c <= 9'b101011010;
				8'b1110000: c <= 9'b110100011;
				8'b1101001: c <= 9'b111100010;
				8'b1110011: c <= 9'b110010;
				8'b1001100: c <= 9'b101101011;
				8'b100001: c <= 9'b101000101;
				8'b1000110: c <= 9'b111001001;
				8'b1110010: c <= 9'b100001001;
				8'b1010000: c <= 9'b111001011;
				8'b1111010: c <= 9'b10010110;
				8'b1010101: c <= 9'b111010100;
				8'b111011: c <= 9'b100010000;
				8'b1001101: c <= 9'b11100101;
				8'b111111: c <= 9'b10;
				8'b1101110: c <= 9'b110101010;
				8'b1111011: c <= 9'b101011;
				8'b1001011: c <= 9'b110110100;
				8'b1101111: c <= 9'b111001100;
				8'b1101000: c <= 9'b1011110;
				8'b101100: c <= 9'b100011011;
				8'b100100: c <= 9'b11001011;
				8'b1111000: c <= 9'b11011100;
				8'b1000101: c <= 9'b11010000;
				8'b1011001: c <= 9'b100000110;
				8'b110100: c <= 9'b110011001;
				8'b1111001: c <= 9'b1111111;
				8'b1110001: c <= 9'b100000001;
				8'b1001111: c <= 9'b1001010;
				8'b1100101: c <= 9'b10111101;
				8'b1111110: c <= 9'b11011101;
				8'b1111100: c <= 9'b100011000;
				8'b1010110: c <= 9'b1011010;
				8'b110010: c <= 9'b111010110;
				8'b1101101: c <= 9'b1101010;
				8'b100011: c <= 9'b111011101;
				8'b1110101: c <= 9'b11001011;
				8'b1111101: c <= 9'b1000110;
				8'b101001: c <= 9'b111100100;
				8'b1010010: c <= 9'b11100101;
				8'b1011000: c <= 9'b101110000;
				8'b101110: c <= 9'b10010011;
				8'b1000001: c <= 9'b100000111;
				default: c <= 9'b0;
			endcase
			9'b110000011 : case(di)
				8'b1000011: c <= 9'b100111111;
				8'b101000: c <= 9'b11001001;
				8'b111010: c <= 9'b11100001;
				8'b110110: c <= 9'b11001111;
				8'b1100100: c <= 9'b110001010;
				8'b1000000: c <= 9'b100110100;
				8'b1110110: c <= 9'b10000111;
				8'b100101: c <= 9'b100110101;
				8'b101111: c <= 9'b10100000;
				8'b100110: c <= 9'b1101000;
				8'b1100011: c <= 9'b1011;
				8'b1001000: c <= 9'b1110011;
				8'b111000: c <= 9'b1110011;
				8'b110001: c <= 9'b110000011;
				8'b1010111: c <= 9'b111110011;
				8'b1001110: c <= 9'b11001010;
				8'b1101010: c <= 9'b101010100;
				8'b1001001: c <= 9'b1111000;
				8'b1100000: c <= 9'b101111110;
				8'b110111: c <= 9'b110100110;
				8'b1011101: c <= 9'b110101001;
				8'b1011011: c <= 9'b11011001;
				8'b111001: c <= 9'b111101110;
				8'b1001010: c <= 9'b100100111;
				8'b110011: c <= 9'b10100010;
				8'b1101100: c <= 9'b110111110;
				8'b1110111: c <= 9'b1011000;
				8'b101011: c <= 9'b110001101;
				8'b1101011: c <= 9'b100101101;
				8'b111100: c <= 9'b101010010;
				8'b1000111: c <= 9'b110011101;
				8'b1011111: c <= 9'b100100010;
				8'b1110100: c <= 9'b101001001;
				8'b101101: c <= 9'b1111010;
				8'b1010011: c <= 9'b1;
				8'b1100001: c <= 9'b10110110;
				8'b110101: c <= 9'b111111101;
				8'b1000100: c <= 9'b111111011;
				8'b1010001: c <= 9'b10111110;
				8'b1010100: c <= 9'b11010;
				8'b1100110: c <= 9'b111001011;
				8'b101010: c <= 9'b101011111;
				8'b1011110: c <= 9'b10100100;
				8'b1100111: c <= 9'b110111000;
				8'b1011010: c <= 9'b101100;
				8'b1000010: c <= 9'b110;
				8'b111101: c <= 9'b101010001;
				8'b110000: c <= 9'b10001110;
				8'b111110: c <= 9'b111001010;
				8'b1100010: c <= 9'b11110001;
				8'b1110000: c <= 9'b101010;
				8'b1101001: c <= 9'b100001101;
				8'b1110011: c <= 9'b11001101;
				8'b1001100: c <= 9'b1010000;
				8'b100001: c <= 9'b101100001;
				8'b1000110: c <= 9'b10110110;
				8'b1110010: c <= 9'b10000;
				8'b1010000: c <= 9'b10110100;
				8'b1111010: c <= 9'b10010110;
				8'b1010101: c <= 9'b10100100;
				8'b111011: c <= 9'b10010101;
				8'b1001101: c <= 9'b100101;
				8'b111111: c <= 9'b110010001;
				8'b1101110: c <= 9'b100011101;
				8'b1111011: c <= 9'b101001110;
				8'b1001011: c <= 9'b11101001;
				8'b1101111: c <= 9'b1000011;
				8'b1101000: c <= 9'b110000000;
				8'b101100: c <= 9'b110101100;
				8'b100100: c <= 9'b1010010;
				8'b1111000: c <= 9'b1110010;
				8'b1000101: c <= 9'b101001100;
				8'b1011001: c <= 9'b111001110;
				8'b110100: c <= 9'b101100;
				8'b1111001: c <= 9'b11100101;
				8'b1110001: c <= 9'b111001001;
				8'b1001111: c <= 9'b110100011;
				8'b1100101: c <= 9'b10001111;
				8'b1111110: c <= 9'b110111001;
				8'b1111100: c <= 9'b10110101;
				8'b1010110: c <= 9'b111001111;
				8'b110010: c <= 9'b11000;
				8'b1101101: c <= 9'b11001;
				8'b100011: c <= 9'b101101100;
				8'b1110101: c <= 9'b1;
				8'b1111101: c <= 9'b111010110;
				8'b101001: c <= 9'b10101000;
				8'b1010010: c <= 9'b101011;
				8'b1011000: c <= 9'b11011100;
				8'b101110: c <= 9'b111010001;
				8'b1000001: c <= 9'b1000010;
				default: c <= 9'b0;
			endcase
			9'b11011 : case(di)
				8'b1000011: c <= 9'b101101110;
				8'b101000: c <= 9'b110000101;
				8'b111010: c <= 9'b100100011;
				8'b110110: c <= 9'b110001101;
				8'b1100100: c <= 9'b100100111;
				8'b1000000: c <= 9'b101101000;
				8'b1110110: c <= 9'b11101100;
				8'b100101: c <= 9'b110001001;
				8'b101111: c <= 9'b101001010;
				8'b100110: c <= 9'b10000110;
				8'b1100011: c <= 9'b101100000;
				8'b1001000: c <= 9'b10010001;
				8'b111000: c <= 9'b111100001;
				8'b110001: c <= 9'b101101101;
				8'b1010111: c <= 9'b101110001;
				8'b1001110: c <= 9'b10010111;
				8'b1101010: c <= 9'b111101100;
				8'b1001001: c <= 9'b111010000;
				8'b1100000: c <= 9'b100100010;
				8'b110111: c <= 9'b110111;
				8'b1011101: c <= 9'b111000;
				8'b1011011: c <= 9'b11100100;
				8'b111001: c <= 9'b1000001;
				8'b1001010: c <= 9'b1000111;
				8'b110011: c <= 9'b100011;
				8'b1101100: c <= 9'b110101111;
				8'b1110111: c <= 9'b10100110;
				8'b101011: c <= 9'b110111110;
				8'b1101011: c <= 9'b111110110;
				8'b111100: c <= 9'b101110100;
				8'b1000111: c <= 9'b101010101;
				8'b1011111: c <= 9'b11001101;
				8'b1110100: c <= 9'b1000001;
				8'b101101: c <= 9'b11011011;
				8'b1010011: c <= 9'b111000111;
				8'b1100001: c <= 9'b101000110;
				8'b110101: c <= 9'b11011001;
				8'b1000100: c <= 9'b101011111;
				8'b1010001: c <= 9'b100010101;
				8'b1010100: c <= 9'b10010111;
				8'b1100110: c <= 9'b100000001;
				8'b101010: c <= 9'b11000010;
				8'b1011110: c <= 9'b100101100;
				8'b1100111: c <= 9'b101100001;
				8'b1011010: c <= 9'b100011101;
				8'b1000010: c <= 9'b110011010;
				8'b111101: c <= 9'b101101011;
				8'b110000: c <= 9'b1011;
				8'b111110: c <= 9'b110111110;
				8'b1100010: c <= 9'b110101101;
				8'b1110000: c <= 9'b11010001;
				8'b1101001: c <= 9'b1001100;
				8'b1110011: c <= 9'b10011100;
				8'b1001100: c <= 9'b11000011;
				8'b100001: c <= 9'b110100011;
				8'b1000110: c <= 9'b111110110;
				8'b1110010: c <= 9'b110111010;
				8'b1010000: c <= 9'b1001011;
				8'b1111010: c <= 9'b111110000;
				8'b1010101: c <= 9'b101010010;
				8'b111011: c <= 9'b10111101;
				8'b1001101: c <= 9'b110111111;
				8'b111111: c <= 9'b1100100;
				8'b1101110: c <= 9'b1000111;
				8'b1111011: c <= 9'b100100101;
				8'b1001011: c <= 9'b111001100;
				8'b1101111: c <= 9'b101010111;
				8'b1101000: c <= 9'b10100101;
				8'b101100: c <= 9'b100111000;
				8'b100100: c <= 9'b101001;
				8'b1111000: c <= 9'b1001011;
				8'b1000101: c <= 9'b110100001;
				8'b1011001: c <= 9'b101101100;
				8'b110100: c <= 9'b1111011;
				8'b1111001: c <= 9'b1110101;
				8'b1110001: c <= 9'b11100100;
				8'b1001111: c <= 9'b1000;
				8'b1100101: c <= 9'b1110000;
				8'b1111110: c <= 9'b11001110;
				8'b1111100: c <= 9'b1001001;
				8'b1010110: c <= 9'b1101;
				8'b110010: c <= 9'b10100110;
				8'b1101101: c <= 9'b10000;
				8'b100011: c <= 9'b1010001;
				8'b1110101: c <= 9'b110000110;
				8'b1111101: c <= 9'b10101111;
				8'b101001: c <= 9'b100000111;
				8'b1010010: c <= 9'b111011101;
				8'b1011000: c <= 9'b110011000;
				8'b101110: c <= 9'b11010100;
				8'b1000001: c <= 9'b1000110;
				default: c <= 9'b0;
			endcase
			9'b10010000 : case(di)
				8'b1000011: c <= 9'b101010101;
				8'b101000: c <= 9'b101011101;
				8'b111010: c <= 9'b11101101;
				8'b110110: c <= 9'b11110110;
				8'b1100100: c <= 9'b110011101;
				8'b1000000: c <= 9'b10011011;
				8'b1110110: c <= 9'b110111011;
				8'b100101: c <= 9'b11101100;
				8'b101111: c <= 9'b10000110;
				8'b100110: c <= 9'b111100111;
				8'b1100011: c <= 9'b111001100;
				8'b1001000: c <= 9'b110000101;
				8'b111000: c <= 9'b1010111;
				8'b110001: c <= 9'b100000110;
				8'b1010111: c <= 9'b110101111;
				8'b1001110: c <= 9'b10100011;
				8'b1101010: c <= 9'b1011011;
				8'b1001001: c <= 9'b10101000;
				8'b1100000: c <= 9'b10110010;
				8'b110111: c <= 9'b1000001;
				8'b1011101: c <= 9'b110111111;
				8'b1011011: c <= 9'b11101001;
				8'b111001: c <= 9'b100110;
				8'b1001010: c <= 9'b10110;
				8'b110011: c <= 9'b110010001;
				8'b1101100: c <= 9'b11110001;
				8'b1110111: c <= 9'b1000101;
				8'b101011: c <= 9'b11111001;
				8'b1101011: c <= 9'b100101;
				8'b111100: c <= 9'b10111111;
				8'b1000111: c <= 9'b1100000;
				8'b1011111: c <= 9'b101000001;
				8'b1110100: c <= 9'b1001101;
				8'b101101: c <= 9'b10001011;
				8'b1010011: c <= 9'b111100001;
				8'b1100001: c <= 9'b101000011;
				8'b110101: c <= 9'b101001;
				8'b1000100: c <= 9'b110101111;
				8'b1010001: c <= 9'b110011010;
				8'b1010100: c <= 9'b11110111;
				8'b1100110: c <= 9'b11110000;
				8'b101010: c <= 9'b11101111;
				8'b1011110: c <= 9'b101010110;
				8'b1100111: c <= 9'b1101000;
				8'b1011010: c <= 9'b110000010;
				8'b1000010: c <= 9'b110110110;
				8'b111101: c <= 9'b100011111;
				8'b110000: c <= 9'b100001011;
				8'b111110: c <= 9'b1000010;
				8'b1100010: c <= 9'b11001000;
				8'b1110000: c <= 9'b10111010;
				8'b1101001: c <= 9'b11011110;
				8'b1110011: c <= 9'b101000011;
				8'b1001100: c <= 9'b101011101;
				8'b100001: c <= 9'b111100110;
				8'b1000110: c <= 9'b111110101;
				8'b1110010: c <= 9'b111110001;
				8'b1010000: c <= 9'b110001010;
				8'b1111010: c <= 9'b100100000;
				8'b1010101: c <= 9'b11110110;
				8'b111011: c <= 9'b101010000;
				8'b1001101: c <= 9'b10001000;
				8'b111111: c <= 9'b111100110;
				8'b1101110: c <= 9'b11100;
				8'b1111011: c <= 9'b101000111;
				8'b1001011: c <= 9'b100011111;
				8'b1101111: c <= 9'b100011000;
				8'b1101000: c <= 9'b110010101;
				8'b101100: c <= 9'b100101101;
				8'b100100: c <= 9'b100101100;
				8'b1111000: c <= 9'b101110101;
				8'b1000101: c <= 9'b10011;
				8'b1011001: c <= 9'b100110010;
				8'b110100: c <= 9'b111001011;
				8'b1111001: c <= 9'b101011010;
				8'b1110001: c <= 9'b11110001;
				8'b1001111: c <= 9'b110111100;
				8'b1100101: c <= 9'b1000110;
				8'b1111110: c <= 9'b10000010;
				8'b1111100: c <= 9'b111001;
				8'b1010110: c <= 9'b11110;
				8'b110010: c <= 9'b11000001;
				8'b1101101: c <= 9'b111000110;
				8'b100011: c <= 9'b110011011;
				8'b1110101: c <= 9'b100001111;
				8'b1111101: c <= 9'b110010100;
				8'b101001: c <= 9'b100110111;
				8'b1010010: c <= 9'b11110100;
				8'b1011000: c <= 9'b1011010;
				8'b101110: c <= 9'b100100111;
				8'b1000001: c <= 9'b111101110;
				default: c <= 9'b0;
			endcase
			9'b101001011 : case(di)
				8'b1000011: c <= 9'b111011100;
				8'b101000: c <= 9'b100010100;
				8'b111010: c <= 9'b11001110;
				8'b110110: c <= 9'b111110110;
				8'b1100100: c <= 9'b110001111;
				8'b1000000: c <= 9'b111011001;
				8'b1110110: c <= 9'b11101111;
				8'b100101: c <= 9'b1000101;
				8'b101111: c <= 9'b10001111;
				8'b100110: c <= 9'b100001011;
				8'b1100011: c <= 9'b111101010;
				8'b1001000: c <= 9'b101000100;
				8'b111000: c <= 9'b10110101;
				8'b110001: c <= 9'b1100100;
				8'b1010111: c <= 9'b110111010;
				8'b1001110: c <= 9'b11011000;
				8'b1101010: c <= 9'b1100001;
				8'b1001001: c <= 9'b100111111;
				8'b1100000: c <= 9'b10010011;
				8'b110111: c <= 9'b100001110;
				8'b1011101: c <= 9'b11001010;
				8'b1011011: c <= 9'b11010101;
				8'b111001: c <= 9'b1000010;
				8'b1001010: c <= 9'b110010;
				8'b110011: c <= 9'b110100101;
				8'b1101100: c <= 9'b10111000;
				8'b1110111: c <= 9'b111011010;
				8'b101011: c <= 9'b11111001;
				8'b1101011: c <= 9'b11001011;
				8'b111100: c <= 9'b10001101;
				8'b1000111: c <= 9'b111010111;
				8'b1011111: c <= 9'b1000010;
				8'b1110100: c <= 9'b111111;
				8'b101101: c <= 9'b111110011;
				8'b1010011: c <= 9'b110001110;
				8'b1100001: c <= 9'b110011010;
				8'b110101: c <= 9'b101110101;
				8'b1000100: c <= 9'b10100011;
				8'b1010001: c <= 9'b100010001;
				8'b1010100: c <= 9'b101001011;
				8'b1100110: c <= 9'b101100110;
				8'b101010: c <= 9'b1001100;
				8'b1011110: c <= 9'b100001;
				8'b1100111: c <= 9'b1001101;
				8'b1011010: c <= 9'b110111010;
				8'b1000010: c <= 9'b100111000;
				8'b111101: c <= 9'b101101101;
				8'b110000: c <= 9'b101000;
				8'b111110: c <= 9'b101110;
				8'b1100010: c <= 9'b110010;
				8'b1110000: c <= 9'b10011100;
				8'b1101001: c <= 9'b10;
				8'b1110011: c <= 9'b11010011;
				8'b1001100: c <= 9'b10001111;
				8'b100001: c <= 9'b100000100;
				8'b1000110: c <= 9'b110011001;
				8'b1110010: c <= 9'b101010000;
				8'b1010000: c <= 9'b101101001;
				8'b1111010: c <= 9'b10010;
				8'b1010101: c <= 9'b11110011;
				8'b111011: c <= 9'b111101100;
				8'b1001101: c <= 9'b100111011;
				8'b111111: c <= 9'b111100101;
				8'b1101110: c <= 9'b111001;
				8'b1111011: c <= 9'b110110;
				8'b1001011: c <= 9'b100101001;
				8'b1101111: c <= 9'b100100010;
				8'b1101000: c <= 9'b111000;
				8'b101100: c <= 9'b110011111;
				8'b100100: c <= 9'b10001101;
				8'b1111000: c <= 9'b111101;
				8'b1000101: c <= 9'b10001100;
				8'b1011001: c <= 9'b100011100;
				8'b110100: c <= 9'b101111010;
				8'b1111001: c <= 9'b10000001;
				8'b1110001: c <= 9'b1000100;
				8'b1001111: c <= 9'b11110001;
				8'b1100101: c <= 9'b11110111;
				8'b1111110: c <= 9'b10001000;
				8'b1111100: c <= 9'b100111110;
				8'b1010110: c <= 9'b100011000;
				8'b110010: c <= 9'b101100000;
				8'b1101101: c <= 9'b101000101;
				8'b100011: c <= 9'b101000;
				8'b1110101: c <= 9'b11010;
				8'b1111101: c <= 9'b111101010;
				8'b101001: c <= 9'b11010000;
				8'b1010010: c <= 9'b11010000;
				8'b1011000: c <= 9'b10101101;
				8'b101110: c <= 9'b110000010;
				8'b1000001: c <= 9'b111100;
				default: c <= 9'b0;
			endcase
			9'b110000001 : case(di)
				8'b1000011: c <= 9'b10010001;
				8'b101000: c <= 9'b111010001;
				8'b111010: c <= 9'b10000000;
				8'b110110: c <= 9'b10101011;
				8'b1100100: c <= 9'b111111;
				8'b1000000: c <= 9'b1001111;
				8'b1110110: c <= 9'b111100100;
				8'b100101: c <= 9'b111100100;
				8'b101111: c <= 9'b110100010;
				8'b100110: c <= 9'b10011101;
				8'b1100011: c <= 9'b10000000;
				8'b1001000: c <= 9'b1100011;
				8'b111000: c <= 9'b111110000;
				8'b110001: c <= 9'b110111;
				8'b1010111: c <= 9'b101001;
				8'b1001110: c <= 9'b110001101;
				8'b1101010: c <= 9'b10110100;
				8'b1001001: c <= 9'b101111010;
				8'b1100000: c <= 9'b10111001;
				8'b110111: c <= 9'b11010111;
				8'b1011101: c <= 9'b101000100;
				8'b1011011: c <= 9'b11101001;
				8'b111001: c <= 9'b10100111;
				8'b1001010: c <= 9'b10101000;
				8'b110011: c <= 9'b11001101;
				8'b1101100: c <= 9'b10101;
				8'b1110111: c <= 9'b1011111;
				8'b101011: c <= 9'b10100110;
				8'b1101011: c <= 9'b111000000;
				8'b111100: c <= 9'b10110001;
				8'b1000111: c <= 9'b10010101;
				8'b1011111: c <= 9'b10111110;
				8'b1110100: c <= 9'b11010111;
				8'b101101: c <= 9'b100000111;
				8'b1010011: c <= 9'b1111010;
				8'b1100001: c <= 9'b111010000;
				8'b110101: c <= 9'b100100;
				8'b1000100: c <= 9'b11001001;
				8'b1010001: c <= 9'b111001010;
				8'b1010100: c <= 9'b1011000;
				8'b1100110: c <= 9'b101110010;
				8'b101010: c <= 9'b101110100;
				8'b1011110: c <= 9'b101001010;
				8'b1100111: c <= 9'b111010010;
				8'b1011010: c <= 9'b10110010;
				8'b1000010: c <= 9'b111110011;
				8'b111101: c <= 9'b1000110;
				8'b110000: c <= 9'b1010001;
				8'b111110: c <= 9'b11000;
				8'b1100010: c <= 9'b11011100;
				8'b1110000: c <= 9'b111110000;
				8'b1101001: c <= 9'b111001111;
				8'b1110011: c <= 9'b111010110;
				8'b1001100: c <= 9'b1110011;
				8'b100001: c <= 9'b110011111;
				8'b1000110: c <= 9'b11111000;
				8'b1110010: c <= 9'b1100011;
				8'b1010000: c <= 9'b110011;
				8'b1111010: c <= 9'b1010001;
				8'b1010101: c <= 9'b100111011;
				8'b111011: c <= 9'b100101;
				8'b1001101: c <= 9'b10001010;
				8'b111111: c <= 9'b110110;
				8'b1101110: c <= 9'b111100010;
				8'b1111011: c <= 9'b110100101;
				8'b1001011: c <= 9'b110100010;
				8'b1101111: c <= 9'b101001111;
				8'b1101000: c <= 9'b111001100;
				8'b101100: c <= 9'b1001011;
				8'b100100: c <= 9'b11111000;
				8'b1111000: c <= 9'b11110110;
				8'b1000101: c <= 9'b101001010;
				8'b1011001: c <= 9'b1011010;
				8'b110100: c <= 9'b100100000;
				8'b1111001: c <= 9'b100001;
				8'b1110001: c <= 9'b100111000;
				8'b1001111: c <= 9'b10111010;
				8'b1100101: c <= 9'b10111101;
				8'b1111110: c <= 9'b110000010;
				8'b1111100: c <= 9'b111010110;
				8'b1010110: c <= 9'b10101101;
				8'b110010: c <= 9'b10000010;
				8'b1101101: c <= 9'b10010000;
				8'b100011: c <= 9'b11110011;
				8'b1110101: c <= 9'b101001000;
				8'b1111101: c <= 9'b1110001;
				8'b101001: c <= 9'b101101110;
				8'b1010010: c <= 9'b10010100;
				8'b1011000: c <= 9'b1111011;
				8'b101110: c <= 9'b1111001;
				8'b1000001: c <= 9'b1100001;
				default: c <= 9'b0;
			endcase
			9'b111111011 : case(di)
				8'b1000011: c <= 9'b10101;
				8'b101000: c <= 9'b110101101;
				8'b111010: c <= 9'b10011101;
				8'b110110: c <= 9'b110000010;
				8'b1100100: c <= 9'b10101101;
				8'b1000000: c <= 9'b101111000;
				8'b1110110: c <= 9'b110001011;
				8'b100101: c <= 9'b111101000;
				8'b101111: c <= 9'b100110111;
				8'b100110: c <= 9'b111011;
				8'b1100011: c <= 9'b1011011;
				8'b1001000: c <= 9'b10000;
				8'b111000: c <= 9'b110000010;
				8'b110001: c <= 9'b1010110;
				8'b1010111: c <= 9'b1111;
				8'b1001110: c <= 9'b110001011;
				8'b1101010: c <= 9'b111000100;
				8'b1001001: c <= 9'b101011101;
				8'b1100000: c <= 9'b111111010;
				8'b110111: c <= 9'b11001000;
				8'b1011101: c <= 9'b111001110;
				8'b1011011: c <= 9'b100100111;
				8'b111001: c <= 9'b1000101;
				8'b1001010: c <= 9'b1100100;
				8'b110011: c <= 9'b100110100;
				8'b1101100: c <= 9'b100111011;
				8'b1110111: c <= 9'b1111101;
				8'b101011: c <= 9'b110011111;
				8'b1101011: c <= 9'b1101100;
				8'b111100: c <= 9'b110100101;
				8'b1000111: c <= 9'b11111010;
				8'b1011111: c <= 9'b11101011;
				8'b1110100: c <= 9'b100010000;
				8'b101101: c <= 9'b110001;
				8'b1010011: c <= 9'b11101000;
				8'b1100001: c <= 9'b10010100;
				8'b110101: c <= 9'b1010101;
				8'b1000100: c <= 9'b1110100;
				8'b1010001: c <= 9'b1001111;
				8'b1010100: c <= 9'b111111101;
				8'b1100110: c <= 9'b11101;
				8'b101010: c <= 9'b100101000;
				8'b1011110: c <= 9'b100001011;
				8'b1100111: c <= 9'b10110110;
				8'b1011010: c <= 9'b10001001;
				8'b1000010: c <= 9'b1100;
				8'b111101: c <= 9'b1101001;
				8'b110000: c <= 9'b100011000;
				8'b111110: c <= 9'b111011;
				8'b1100010: c <= 9'b101001000;
				8'b1110000: c <= 9'b110101100;
				8'b1101001: c <= 9'b101110011;
				8'b1110011: c <= 9'b101100;
				8'b1001100: c <= 9'b111000011;
				8'b100001: c <= 9'b110111111;
				8'b1000110: c <= 9'b1011110;
				8'b1110010: c <= 9'b11011011;
				8'b1010000: c <= 9'b10001100;
				8'b1111010: c <= 9'b1011110;
				8'b1010101: c <= 9'b110011111;
				8'b111011: c <= 9'b101110010;
				8'b1001101: c <= 9'b11001010;
				8'b111111: c <= 9'b1111110;
				8'b1101110: c <= 9'b100100010;
				8'b1111011: c <= 9'b10110111;
				8'b1001011: c <= 9'b111010110;
				8'b1101111: c <= 9'b101100111;
				8'b1101000: c <= 9'b11110011;
				8'b101100: c <= 9'b10100110;
				8'b100100: c <= 9'b110100100;
				8'b1111000: c <= 9'b1010110;
				8'b1000101: c <= 9'b100110011;
				8'b1011001: c <= 9'b100100000;
				8'b110100: c <= 9'b101010110;
				8'b1111001: c <= 9'b10100000;
				8'b1110001: c <= 9'b100001110;
				8'b1001111: c <= 9'b101101011;
				8'b1100101: c <= 9'b11;
				8'b1111110: c <= 9'b10110111;
				8'b1111100: c <= 9'b101000010;
				8'b1010110: c <= 9'b1100000;
				8'b110010: c <= 9'b100010111;
				8'b1101101: c <= 9'b10001101;
				8'b100011: c <= 9'b11101000;
				8'b1110101: c <= 9'b110101011;
				8'b1111101: c <= 9'b10010001;
				8'b101001: c <= 9'b1001011;
				8'b1010010: c <= 9'b110011;
				8'b1011000: c <= 9'b1011010;
				8'b101110: c <= 9'b1111000;
				8'b1000001: c <= 9'b101110010;
				default: c <= 9'b0;
			endcase
			9'b10000011 : case(di)
				8'b1000011: c <= 9'b101010;
				8'b101000: c <= 9'b111100000;
				8'b111010: c <= 9'b10100100;
				8'b110110: c <= 9'b110010010;
				8'b1100100: c <= 9'b10011000;
				8'b1000000: c <= 9'b101001;
				8'b1110110: c <= 9'b111100111;
				8'b100101: c <= 9'b111111000;
				8'b101111: c <= 9'b101001001;
				8'b100110: c <= 9'b100001010;
				8'b1100011: c <= 9'b11001000;
				8'b1001000: c <= 9'b100110100;
				8'b111000: c <= 9'b100000100;
				8'b110001: c <= 9'b101100110;
				8'b1010111: c <= 9'b110010;
				8'b1001110: c <= 9'b11000011;
				8'b1101010: c <= 9'b100011;
				8'b1001001: c <= 9'b100001010;
				8'b1100000: c <= 9'b1;
				8'b110111: c <= 9'b111111101;
				8'b1011101: c <= 9'b110001;
				8'b1011011: c <= 9'b110111010;
				8'b111001: c <= 9'b110100000;
				8'b1001010: c <= 9'b110101011;
				8'b110011: c <= 9'b111011001;
				8'b1101100: c <= 9'b10110111;
				8'b1110111: c <= 9'b1101010;
				8'b101011: c <= 9'b100110101;
				8'b1101011: c <= 9'b111101101;
				8'b111100: c <= 9'b11100001;
				8'b1000111: c <= 9'b11010010;
				8'b1011111: c <= 9'b10100110;
				8'b1110100: c <= 9'b101010101;
				8'b101101: c <= 9'b101;
				8'b1010011: c <= 9'b110111011;
				8'b1100001: c <= 9'b1011111;
				8'b110101: c <= 9'b110111110;
				8'b1000100: c <= 9'b10101;
				8'b1010001: c <= 9'b10110111;
				8'b1010100: c <= 9'b111010100;
				8'b1100110: c <= 9'b111101111;
				8'b101010: c <= 9'b11011101;
				8'b1011110: c <= 9'b10010011;
				8'b1100111: c <= 9'b110001111;
				8'b1011010: c <= 9'b111111;
				8'b1000010: c <= 9'b110000010;
				8'b111101: c <= 9'b110111100;
				8'b110000: c <= 9'b111101101;
				8'b111110: c <= 9'b10001001;
				8'b1100010: c <= 9'b100001110;
				8'b1110000: c <= 9'b1011001;
				8'b1101001: c <= 9'b10011100;
				8'b1110011: c <= 9'b11111;
				8'b1001100: c <= 9'b1100010;
				8'b100001: c <= 9'b10111101;
				8'b1000110: c <= 9'b111101;
				8'b1110010: c <= 9'b100001011;
				8'b1010000: c <= 9'b100101110;
				8'b1111010: c <= 9'b110010111;
				8'b1010101: c <= 9'b11101000;
				8'b111011: c <= 9'b110111010;
				8'b1001101: c <= 9'b1001011;
				8'b111111: c <= 9'b110011001;
				8'b1101110: c <= 9'b111101101;
				8'b1111011: c <= 9'b100101100;
				8'b1001011: c <= 9'b101000011;
				8'b1101111: c <= 9'b10101001;
				8'b1101000: c <= 9'b100001110;
				8'b101100: c <= 9'b1111101;
				8'b100100: c <= 9'b101111001;
				8'b1111000: c <= 9'b11100011;
				8'b1000101: c <= 9'b10010111;
				8'b1011001: c <= 9'b10;
				8'b110100: c <= 9'b110011001;
				8'b1111001: c <= 9'b11010100;
				8'b1110001: c <= 9'b110111100;
				8'b1001111: c <= 9'b100010110;
				8'b1100101: c <= 9'b10;
				8'b1111110: c <= 9'b10010110;
				8'b1111100: c <= 9'b110001111;
				8'b1010110: c <= 9'b110100001;
				8'b110010: c <= 9'b110101100;
				8'b1101101: c <= 9'b10011;
				8'b100011: c <= 9'b10101110;
				8'b1110101: c <= 9'b111111000;
				8'b1111101: c <= 9'b111011001;
				8'b101001: c <= 9'b10100;
				8'b1010010: c <= 9'b100101110;
				8'b1011000: c <= 9'b11101000;
				8'b101110: c <= 9'b101110110;
				8'b1000001: c <= 9'b11101011;
				default: c <= 9'b0;
			endcase
			9'b1101101 : case(di)
				8'b1000011: c <= 9'b100;
				8'b101000: c <= 9'b111011;
				8'b111010: c <= 9'b11100100;
				8'b110110: c <= 9'b10001000;
				8'b1100100: c <= 9'b11111010;
				8'b1000000: c <= 9'b100001110;
				8'b1110110: c <= 9'b1110011;
				8'b100101: c <= 9'b1000100;
				8'b101111: c <= 9'b1111001;
				8'b100110: c <= 9'b1110100;
				8'b1100011: c <= 9'b10010011;
				8'b1001000: c <= 9'b10000010;
				8'b111000: c <= 9'b10011010;
				8'b110001: c <= 9'b11001000;
				8'b1010111: c <= 9'b111001011;
				8'b1001110: c <= 9'b100101;
				8'b1101010: c <= 9'b10110010;
				8'b1001001: c <= 9'b101001011;
				8'b1100000: c <= 9'b111111110;
				8'b110111: c <= 9'b100000010;
				8'b1011101: c <= 9'b111001001;
				8'b1011011: c <= 9'b111101010;
				8'b111001: c <= 9'b10111101;
				8'b1001010: c <= 9'b110011010;
				8'b110011: c <= 9'b11110101;
				8'b1101100: c <= 9'b100010;
				8'b1110111: c <= 9'b101100111;
				8'b101011: c <= 9'b101001110;
				8'b1101011: c <= 9'b110010011;
				8'b111100: c <= 9'b110100001;
				8'b1000111: c <= 9'b1111010;
				8'b1011111: c <= 9'b10000101;
				8'b1110100: c <= 9'b11111011;
				8'b101101: c <= 9'b11010000;
				8'b1010011: c <= 9'b10101001;
				8'b1100001: c <= 9'b101101111;
				8'b110101: c <= 9'b1110101;
				8'b1000100: c <= 9'b101011001;
				8'b1010001: c <= 9'b1101110;
				8'b1010100: c <= 9'b100101101;
				8'b1100110: c <= 9'b1001100;
				8'b101010: c <= 9'b1000000;
				8'b1011110: c <= 9'b110110000;
				8'b1100111: c <= 9'b110101011;
				8'b1011010: c <= 9'b111010001;
				8'b1000010: c <= 9'b10001001;
				8'b111101: c <= 9'b101111000;
				8'b110000: c <= 9'b1001111;
				8'b111110: c <= 9'b1101000;
				8'b1100010: c <= 9'b100000000;
				8'b1110000: c <= 9'b10111001;
				8'b1101001: c <= 9'b1001;
				8'b1110011: c <= 9'b10010110;
				8'b1001100: c <= 9'b10111;
				8'b100001: c <= 9'b110111001;
				8'b1000110: c <= 9'b101101111;
				8'b1110010: c <= 9'b110100001;
				8'b1010000: c <= 9'b11011010;
				8'b1111010: c <= 9'b11011101;
				8'b1010101: c <= 9'b101010011;
				8'b111011: c <= 9'b101111001;
				8'b1001101: c <= 9'b100101100;
				8'b111111: c <= 9'b101001110;
				8'b1101110: c <= 9'b1000001;
				8'b1111011: c <= 9'b11001;
				8'b1001011: c <= 9'b101100;
				8'b1101111: c <= 9'b100010011;
				8'b1101000: c <= 9'b11111110;
				8'b101100: c <= 9'b100110100;
				8'b100100: c <= 9'b110111110;
				8'b1111000: c <= 9'b110010100;
				8'b1000101: c <= 9'b110111100;
				8'b1011001: c <= 9'b10011000;
				8'b110100: c <= 9'b10110010;
				8'b1111001: c <= 9'b100000110;
				8'b1110001: c <= 9'b1011110;
				8'b1001111: c <= 9'b111100010;
				8'b1100101: c <= 9'b111001110;
				8'b1111110: c <= 9'b1001110;
				8'b1111100: c <= 9'b101011111;
				8'b1010110: c <= 9'b100101111;
				8'b110010: c <= 9'b11110010;
				8'b1101101: c <= 9'b101110001;
				8'b100011: c <= 9'b111111101;
				8'b1110101: c <= 9'b101010000;
				8'b1111101: c <= 9'b111000;
				8'b101001: c <= 9'b101001011;
				8'b1010010: c <= 9'b101001111;
				8'b1011000: c <= 9'b11100110;
				8'b101110: c <= 9'b10;
				8'b1000001: c <= 9'b1;
				default: c <= 9'b0;
			endcase
			9'b11101011 : case(di)
				8'b1000011: c <= 9'b110100110;
				8'b101000: c <= 9'b111110110;
				8'b111010: c <= 9'b1101100;
				8'b110110: c <= 9'b101111111;
				8'b1100100: c <= 9'b100101;
				8'b1000000: c <= 9'b110001001;
				8'b1110110: c <= 9'b110011101;
				8'b100101: c <= 9'b10000101;
				8'b101111: c <= 9'b11011;
				8'b100110: c <= 9'b10000011;
				8'b1100011: c <= 9'b100110000;
				8'b1001000: c <= 9'b1111010;
				8'b111000: c <= 9'b110110010;
				8'b110001: c <= 9'b11001100;
				8'b1010111: c <= 9'b101011000;
				8'b1001110: c <= 9'b111100011;
				8'b1101010: c <= 9'b111000010;
				8'b1001001: c <= 9'b1010011;
				8'b1100000: c <= 9'b10111100;
				8'b110111: c <= 9'b101001110;
				8'b1011101: c <= 9'b100000011;
				8'b1011011: c <= 9'b11011011;
				8'b111001: c <= 9'b10011000;
				8'b1001010: c <= 9'b110011110;
				8'b110011: c <= 9'b100011001;
				8'b1101100: c <= 9'b101011;
				8'b1110111: c <= 9'b101010000;
				8'b101011: c <= 9'b101111001;
				8'b1101011: c <= 9'b110100001;
				8'b111100: c <= 9'b11001000;
				8'b1000111: c <= 9'b10010000;
				8'b1011111: c <= 9'b10110110;
				8'b1110100: c <= 9'b110100011;
				8'b101101: c <= 9'b101100;
				8'b1010011: c <= 9'b11100110;
				8'b1100001: c <= 9'b11101111;
				8'b110101: c <= 9'b10010110;
				8'b1000100: c <= 9'b1100001;
				8'b1010001: c <= 9'b11011010;
				8'b1010100: c <= 9'b100000101;
				8'b1100110: c <= 9'b1101;
				8'b101010: c <= 9'b110001101;
				8'b1011110: c <= 9'b110001100;
				8'b1100111: c <= 9'b10101010;
				8'b1011010: c <= 9'b11101011;
				8'b1000010: c <= 9'b101000001;
				8'b111101: c <= 9'b1110001;
				8'b110000: c <= 9'b101100;
				8'b111110: c <= 9'b10001110;
				8'b1100010: c <= 9'b11110011;
				8'b1110000: c <= 9'b100011;
				8'b1101001: c <= 9'b1011;
				8'b1110011: c <= 9'b11111101;
				8'b1001100: c <= 9'b11111101;
				8'b100001: c <= 9'b101001010;
				8'b1000110: c <= 9'b100001110;
				8'b1110010: c <= 9'b101010011;
				8'b1010000: c <= 9'b101011011;
				8'b1111010: c <= 9'b100101111;
				8'b1010101: c <= 9'b100111111;
				8'b111011: c <= 9'b11000001;
				8'b1001101: c <= 9'b10001100;
				8'b111111: c <= 9'b11000000;
				8'b1101110: c <= 9'b101010;
				8'b1111011: c <= 9'b10010101;
				8'b1001011: c <= 9'b11010100;
				8'b1101111: c <= 9'b100001010;
				8'b1101000: c <= 9'b100100110;
				8'b101100: c <= 9'b111101000;
				8'b100100: c <= 9'b101;
				8'b1111000: c <= 9'b11110111;
				8'b1000101: c <= 9'b101;
				8'b1011001: c <= 9'b100101101;
				8'b110100: c <= 9'b10;
				8'b1111001: c <= 9'b110100001;
				8'b1110001: c <= 9'b111011;
				8'b1001111: c <= 9'b11000001;
				8'b1100101: c <= 9'b110010010;
				8'b1111110: c <= 9'b100010111;
				8'b1111100: c <= 9'b110100000;
				8'b1010110: c <= 9'b1101000;
				8'b110010: c <= 9'b100000110;
				8'b1101101: c <= 9'b1010110;
				8'b100011: c <= 9'b110000111;
				8'b1110101: c <= 9'b110110111;
				8'b1111101: c <= 9'b10100100;
				8'b101001: c <= 9'b100011011;
				8'b1010010: c <= 9'b110100111;
				8'b1011000: c <= 9'b111111000;
				8'b101110: c <= 9'b11010011;
				8'b1000001: c <= 9'b1110111;
				default: c <= 9'b0;
			endcase
			9'b10111001 : case(di)
				8'b1000011: c <= 9'b101100010;
				8'b101000: c <= 9'b110001011;
				8'b111010: c <= 9'b110000;
				8'b110110: c <= 9'b11110111;
				8'b1100100: c <= 9'b111111;
				8'b1000000: c <= 9'b100100000;
				8'b1110110: c <= 9'b11001011;
				8'b100101: c <= 9'b110000001;
				8'b101111: c <= 9'b100110110;
				8'b100110: c <= 9'b110111;
				8'b1100011: c <= 9'b101000;
				8'b1001000: c <= 9'b1001001;
				8'b111000: c <= 9'b101100;
				8'b110001: c <= 9'b11111100;
				8'b1010111: c <= 9'b100101010;
				8'b1001110: c <= 9'b10110100;
				8'b1101010: c <= 9'b101100001;
				8'b1001001: c <= 9'b10001001;
				8'b1100000: c <= 9'b110000110;
				8'b110111: c <= 9'b11010100;
				8'b1011101: c <= 9'b110100;
				8'b1011011: c <= 9'b100101011;
				8'b111001: c <= 9'b10010101;
				8'b1001010: c <= 9'b10101000;
				8'b110011: c <= 9'b110100011;
				8'b1101100: c <= 9'b111100011;
				8'b1110111: c <= 9'b111101110;
				8'b101011: c <= 9'b110101110;
				8'b1101011: c <= 9'b1110100;
				8'b111100: c <= 9'b101001000;
				8'b1000111: c <= 9'b110001;
				8'b1011111: c <= 9'b11110100;
				8'b1110100: c <= 9'b101100010;
				8'b101101: c <= 9'b1000010;
				8'b1010011: c <= 9'b1100111;
				8'b1100001: c <= 9'b1000111;
				8'b110101: c <= 9'b101110;
				8'b1000100: c <= 9'b10001001;
				8'b1010001: c <= 9'b10010011;
				8'b1010100: c <= 9'b100010010;
				8'b1100110: c <= 9'b111001101;
				8'b101010: c <= 9'b110100101;
				8'b1011110: c <= 9'b100111010;
				8'b1100111: c <= 9'b110101001;
				8'b1011010: c <= 9'b101001;
				8'b1000010: c <= 9'b10101;
				8'b111101: c <= 9'b101110110;
				8'b110000: c <= 9'b111011010;
				8'b111110: c <= 9'b101010011;
				8'b1100010: c <= 9'b11010101;
				8'b1110000: c <= 9'b11110;
				8'b1101001: c <= 9'b111110001;
				8'b1110011: c <= 9'b1001101;
				8'b1001100: c <= 9'b1101111;
				8'b100001: c <= 9'b10000011;
				8'b1000110: c <= 9'b110001110;
				8'b1110010: c <= 9'b110101;
				8'b1010000: c <= 9'b101010111;
				8'b1111010: c <= 9'b11100010;
				8'b1010101: c <= 9'b111100111;
				8'b111011: c <= 9'b1111011;
				8'b1001101: c <= 9'b10101;
				8'b111111: c <= 9'b101110111;
				8'b1101110: c <= 9'b100010110;
				8'b1111011: c <= 9'b100001001;
				8'b1001011: c <= 9'b1100101;
				8'b1101111: c <= 9'b10110;
				8'b1101000: c <= 9'b11000111;
				8'b101100: c <= 9'b10110011;
				8'b100100: c <= 9'b11100111;
				8'b1111000: c <= 9'b110111010;
				8'b1000101: c <= 9'b101011;
				8'b1011001: c <= 9'b1000101;
				8'b110100: c <= 9'b10001110;
				8'b1111001: c <= 9'b110001;
				8'b1110001: c <= 9'b1011110;
				8'b1001111: c <= 9'b100010001;
				8'b1100101: c <= 9'b11101001;
				8'b1111110: c <= 9'b101100010;
				8'b1111100: c <= 9'b11100100;
				8'b1010110: c <= 9'b101111110;
				8'b110010: c <= 9'b101000001;
				8'b1101101: c <= 9'b10111011;
				8'b100011: c <= 9'b11011;
				8'b1110101: c <= 9'b111010100;
				8'b1111101: c <= 9'b10111111;
				8'b101001: c <= 9'b111001101;
				8'b1010010: c <= 9'b1011000;
				8'b1011000: c <= 9'b10110011;
				8'b101110: c <= 9'b101000101;
				8'b1000001: c <= 9'b11001100;
				default: c <= 9'b0;
			endcase
			9'b101101101 : case(di)
				8'b1000011: c <= 9'b100000011;
				8'b101000: c <= 9'b101001000;
				8'b111010: c <= 9'b11111011;
				8'b110110: c <= 9'b111111;
				8'b1100100: c <= 9'b11010;
				8'b1000000: c <= 9'b10101;
				8'b1110110: c <= 9'b11010000;
				8'b100101: c <= 9'b101100110;
				8'b101111: c <= 9'b10100;
				8'b100110: c <= 9'b101000010;
				8'b1100011: c <= 9'b111010111;
				8'b1001000: c <= 9'b100111100;
				8'b111000: c <= 9'b11010100;
				8'b110001: c <= 9'b100;
				8'b1010111: c <= 9'b101011101;
				8'b1001110: c <= 9'b1100110;
				8'b1101010: c <= 9'b101010010;
				8'b1001001: c <= 9'b100100000;
				8'b1100000: c <= 9'b111101100;
				8'b110111: c <= 9'b111110011;
				8'b1011101: c <= 9'b1111110;
				8'b1011011: c <= 9'b11001100;
				8'b111001: c <= 9'b100111011;
				8'b1001010: c <= 9'b111001101;
				8'b110011: c <= 9'b101001111;
				8'b1101100: c <= 9'b10010011;
				8'b1110111: c <= 9'b1101000;
				8'b101011: c <= 9'b100101111;
				8'b1101011: c <= 9'b101110111;
				8'b111100: c <= 9'b11100001;
				8'b1000111: c <= 9'b1110010;
				8'b1011111: c <= 9'b111111111;
				8'b1110100: c <= 9'b11101011;
				8'b101101: c <= 9'b111100000;
				8'b1010011: c <= 9'b10001000;
				8'b1100001: c <= 9'b10101100;
				8'b110101: c <= 9'b11110001;
				8'b1000100: c <= 9'b1110111;
				8'b1010001: c <= 9'b111111011;
				8'b1010100: c <= 9'b110110010;
				8'b1100110: c <= 9'b1110011;
				8'b101010: c <= 9'b10001010;
				8'b1011110: c <= 9'b1001000;
				8'b1100111: c <= 9'b111101000;
				8'b1011010: c <= 9'b11000011;
				8'b1000010: c <= 9'b10111010;
				8'b111101: c <= 9'b11111;
				8'b110000: c <= 9'b110111;
				8'b111110: c <= 9'b101101110;
				8'b1100010: c <= 9'b100111;
				8'b1110000: c <= 9'b1111111;
				8'b1101001: c <= 9'b10100101;
				8'b1110011: c <= 9'b10100011;
				8'b1001100: c <= 9'b111011010;
				8'b100001: c <= 9'b1011000;
				8'b1000110: c <= 9'b10101011;
				8'b1110010: c <= 9'b101101011;
				8'b1010000: c <= 9'b110100110;
				8'b1111010: c <= 9'b10111001;
				8'b1010101: c <= 9'b100011001;
				8'b111011: c <= 9'b100011001;
				8'b1001101: c <= 9'b11111011;
				8'b111111: c <= 9'b11110000;
				8'b1101110: c <= 9'b10110101;
				8'b1111011: c <= 9'b100111010;
				8'b1001011: c <= 9'b101000001;
				8'b1101111: c <= 9'b111;
				8'b1101000: c <= 9'b1111001;
				8'b101100: c <= 9'b11100101;
				8'b100100: c <= 9'b101001110;
				8'b1111000: c <= 9'b1111110;
				8'b1000101: c <= 9'b101110011;
				8'b1011001: c <= 9'b100011010;
				8'b110100: c <= 9'b100000111;
				8'b1111001: c <= 9'b11101000;
				8'b1110001: c <= 9'b100101101;
				8'b1001111: c <= 9'b10100;
				8'b1100101: c <= 9'b110110100;
				8'b1111110: c <= 9'b111111101;
				8'b1111100: c <= 9'b1001;
				8'b1010110: c <= 9'b10000101;
				8'b110010: c <= 9'b1110101;
				8'b1101101: c <= 9'b1111011;
				8'b100011: c <= 9'b1100000;
				8'b1110101: c <= 9'b100000000;
				8'b1111101: c <= 9'b1001011;
				8'b101001: c <= 9'b101011011;
				8'b1010010: c <= 9'b10010011;
				8'b1011000: c <= 9'b1101010;
				8'b101110: c <= 9'b11110110;
				8'b1000001: c <= 9'b101101000;
				default: c <= 9'b0;
			endcase
			9'b110001000 : case(di)
				8'b1000011: c <= 9'b101100;
				8'b101000: c <= 9'b11111011;
				8'b111010: c <= 9'b100110011;
				8'b110110: c <= 9'b111011011;
				8'b1100100: c <= 9'b111111010;
				8'b1000000: c <= 9'b101111000;
				8'b1110110: c <= 9'b11011011;
				8'b100101: c <= 9'b11000000;
				8'b101111: c <= 9'b1101111;
				8'b100110: c <= 9'b101000011;
				8'b1100011: c <= 9'b1110101;
				8'b1001000: c <= 9'b101011011;
				8'b111000: c <= 9'b1100;
				8'b110001: c <= 9'b11010100;
				8'b1010111: c <= 9'b110011100;
				8'b1001110: c <= 9'b101000111;
				8'b1101010: c <= 9'b111101010;
				8'b1001001: c <= 9'b10100100;
				8'b1100000: c <= 9'b10010110;
				8'b110111: c <= 9'b11110;
				8'b1011101: c <= 9'b110100001;
				8'b1011011: c <= 9'b100010110;
				8'b111001: c <= 9'b10101010;
				8'b1001010: c <= 9'b1111011;
				8'b110011: c <= 9'b10111100;
				8'b1101100: c <= 9'b100011011;
				8'b1110111: c <= 9'b101010110;
				8'b101011: c <= 9'b111100;
				8'b1101011: c <= 9'b111100101;
				8'b111100: c <= 9'b101100111;
				8'b1000111: c <= 9'b110001001;
				8'b1011111: c <= 9'b100011;
				8'b1110100: c <= 9'b110000;
				8'b101101: c <= 9'b11010011;
				8'b1010011: c <= 9'b111001110;
				8'b1100001: c <= 9'b100001110;
				8'b110101: c <= 9'b111011110;
				8'b1000100: c <= 9'b11100111;
				8'b1010001: c <= 9'b111100011;
				8'b1010100: c <= 9'b111100;
				8'b1100110: c <= 9'b110111;
				8'b101010: c <= 9'b10001010;
				8'b1011110: c <= 9'b10101100;
				8'b1100111: c <= 9'b10111;
				8'b1011010: c <= 9'b101011001;
				8'b1000010: c <= 9'b1111000;
				8'b111101: c <= 9'b10010011;
				8'b110000: c <= 9'b11110101;
				8'b111110: c <= 9'b100001100;
				8'b1100010: c <= 9'b100001001;
				8'b1110000: c <= 9'b110100100;
				8'b1101001: c <= 9'b100111010;
				8'b1110011: c <= 9'b10001010;
				8'b1001100: c <= 9'b11110;
				8'b100001: c <= 9'b101011001;
				8'b1000110: c <= 9'b1101111;
				8'b1110010: c <= 9'b11001000;
				8'b1010000: c <= 9'b110011;
				8'b1111010: c <= 9'b101111110;
				8'b1010101: c <= 9'b101100;
				8'b111011: c <= 9'b101000001;
				8'b1001101: c <= 9'b10101111;
				8'b111111: c <= 9'b111010;
				8'b1101110: c <= 9'b11111;
				8'b1111011: c <= 9'b11101100;
				8'b1001011: c <= 9'b11011;
				8'b1101111: c <= 9'b10110111;
				8'b1101000: c <= 9'b11110100;
				8'b101100: c <= 9'b111001110;
				8'b100100: c <= 9'b10110101;
				8'b1111000: c <= 9'b111011110;
				8'b1000101: c <= 9'b111110000;
				8'b1011001: c <= 9'b1100001;
				8'b110100: c <= 9'b111100000;
				8'b1111001: c <= 9'b1110011;
				8'b1110001: c <= 9'b11100111;
				8'b1001111: c <= 9'b100111111;
				8'b1100101: c <= 9'b101100000;
				8'b1111110: c <= 9'b101011110;
				8'b1111100: c <= 9'b11010;
				8'b1010110: c <= 9'b100100101;
				8'b110010: c <= 9'b101011111;
				8'b1101101: c <= 9'b110101101;
				8'b100011: c <= 9'b10100111;
				8'b1110101: c <= 9'b100000010;
				8'b1111101: c <= 9'b100011101;
				8'b101001: c <= 9'b111010010;
				8'b1010010: c <= 9'b1111;
				8'b1011000: c <= 9'b111011001;
				8'b101110: c <= 9'b11011100;
				8'b1000001: c <= 9'b1100101;
				default: c <= 9'b0;
			endcase
			9'b111101100 : case(di)
				8'b1000011: c <= 9'b111101010;
				8'b101000: c <= 9'b100111101;
				8'b111010: c <= 9'b101100000;
				8'b110110: c <= 9'b11011011;
				8'b1100100: c <= 9'b1110;
				8'b1000000: c <= 9'b1110;
				8'b1110110: c <= 9'b101110001;
				8'b100101: c <= 9'b11111000;
				8'b101111: c <= 9'b10010111;
				8'b100110: c <= 9'b110011001;
				8'b1100011: c <= 9'b11110111;
				8'b1001000: c <= 9'b11100110;
				8'b111000: c <= 9'b11000010;
				8'b110001: c <= 9'b101110010;
				8'b1010111: c <= 9'b101001;
				8'b1001110: c <= 9'b101101;
				8'b1101010: c <= 9'b111111000;
				8'b1001001: c <= 9'b10000000;
				8'b1100000: c <= 9'b100000110;
				8'b110111: c <= 9'b111111;
				8'b1011101: c <= 9'b1001101;
				8'b1011011: c <= 9'b111011101;
				8'b111001: c <= 9'b11110010;
				8'b1001010: c <= 9'b1100001;
				8'b110011: c <= 9'b10101111;
				8'b1101100: c <= 9'b101000110;
				8'b1110111: c <= 9'b10111001;
				8'b101011: c <= 9'b111001000;
				8'b1101011: c <= 9'b100100110;
				8'b111100: c <= 9'b100001001;
				8'b1000111: c <= 9'b101111110;
				8'b1011111: c <= 9'b10001100;
				8'b1110100: c <= 9'b1;
				8'b101101: c <= 9'b11001010;
				8'b1010011: c <= 9'b10001110;
				8'b1100001: c <= 9'b1111010;
				8'b110101: c <= 9'b11011010;
				8'b1000100: c <= 9'b10100011;
				8'b1010001: c <= 9'b11100010;
				8'b1010100: c <= 9'b110011101;
				8'b1100110: c <= 9'b11001100;
				8'b101010: c <= 9'b101010111;
				8'b1011110: c <= 9'b100000101;
				8'b1100111: c <= 9'b11101011;
				8'b1011010: c <= 9'b10011;
				8'b1000010: c <= 9'b1110010;
				8'b111101: c <= 9'b110100010;
				8'b110000: c <= 9'b1111111;
				8'b111110: c <= 9'b10111100;
				8'b1100010: c <= 9'b101100;
				8'b1110000: c <= 9'b101010101;
				8'b1101001: c <= 9'b110110010;
				8'b1110011: c <= 9'b110010100;
				8'b1001100: c <= 9'b111001100;
				8'b100001: c <= 9'b110001101;
				8'b1000110: c <= 9'b10111110;
				8'b1110010: c <= 9'b1000111;
				8'b1010000: c <= 9'b1001110;
				8'b1111010: c <= 9'b10011111;
				8'b1010101: c <= 9'b11111101;
				8'b111011: c <= 9'b1101110;
				8'b1001101: c <= 9'b11000100;
				8'b111111: c <= 9'b10101101;
				8'b1101110: c <= 9'b110001111;
				8'b1111011: c <= 9'b10100110;
				8'b1001011: c <= 9'b110011101;
				8'b1101111: c <= 9'b10010001;
				8'b1101000: c <= 9'b100111111;
				8'b101100: c <= 9'b1;
				8'b100100: c <= 9'b10000;
				8'b1111000: c <= 9'b1000011;
				8'b1000101: c <= 9'b111001111;
				8'b1011001: c <= 9'b100110111;
				8'b110100: c <= 9'b100101001;
				8'b1111001: c <= 9'b110100011;
				8'b1110001: c <= 9'b111111001;
				8'b1001111: c <= 9'b100100111;
				8'b1100101: c <= 9'b111001001;
				8'b1111110: c <= 9'b1000010;
				8'b1111100: c <= 9'b10011111;
				8'b1010110: c <= 9'b101100111;
				8'b110010: c <= 9'b101100101;
				8'b1101101: c <= 9'b110001110;
				8'b100011: c <= 9'b110010111;
				8'b1110101: c <= 9'b11011001;
				8'b1111101: c <= 9'b10000011;
				8'b101001: c <= 9'b10100000;
				8'b1010010: c <= 9'b110011010;
				8'b1011000: c <= 9'b10001100;
				8'b101110: c <= 9'b100111;
				8'b1000001: c <= 9'b11101001;
				default: c <= 9'b0;
			endcase
			9'b101 : case(di)
				8'b1000011: c <= 9'b10101111;
				8'b101000: c <= 9'b100010010;
				8'b111010: c <= 9'b111100111;
				8'b110110: c <= 9'b110010011;
				8'b1100100: c <= 9'b101000011;
				8'b1000000: c <= 9'b10011101;
				8'b1110110: c <= 9'b110011;
				8'b100101: c <= 9'b101010100;
				8'b101111: c <= 9'b100010101;
				8'b100110: c <= 9'b101111111;
				8'b1100011: c <= 9'b10110010;
				8'b1001000: c <= 9'b1001101;
				8'b111000: c <= 9'b111101111;
				8'b110001: c <= 9'b101111000;
				8'b1010111: c <= 9'b110001000;
				8'b1001110: c <= 9'b111001000;
				8'b1101010: c <= 9'b1010101;
				8'b1001001: c <= 9'b10001010;
				8'b1100000: c <= 9'b110000110;
				8'b110111: c <= 9'b100100;
				8'b1011101: c <= 9'b101111110;
				8'b1011011: c <= 9'b11101100;
				8'b111001: c <= 9'b11011001;
				8'b1001010: c <= 9'b11100110;
				8'b110011: c <= 9'b11100000;
				8'b1101100: c <= 9'b101001000;
				8'b1110111: c <= 9'b110110100;
				8'b101011: c <= 9'b111000101;
				8'b1101011: c <= 9'b110001;
				8'b111100: c <= 9'b110111110;
				8'b1000111: c <= 9'b111101010;
				8'b1011111: c <= 9'b111001011;
				8'b1110100: c <= 9'b110011110;
				8'b101101: c <= 9'b100111110;
				8'b1010011: c <= 9'b11001010;
				8'b1100001: c <= 9'b100101000;
				8'b110101: c <= 9'b111000011;
				8'b1000100: c <= 9'b110111110;
				8'b1010001: c <= 9'b1011111;
				8'b1010100: c <= 9'b10110101;
				8'b1100110: c <= 9'b110110000;
				8'b101010: c <= 9'b111100010;
				8'b1011110: c <= 9'b100010100;
				8'b1100111: c <= 9'b100110000;
				8'b1011010: c <= 9'b101100001;
				8'b1000010: c <= 9'b100100001;
				8'b111101: c <= 9'b10100100;
				8'b110000: c <= 9'b1111100;
				8'b111110: c <= 9'b111111000;
				8'b1100010: c <= 9'b100011001;
				8'b1110000: c <= 9'b110101011;
				8'b1101001: c <= 9'b100100;
				8'b1110011: c <= 9'b110110111;
				8'b1001100: c <= 9'b111010110;
				8'b100001: c <= 9'b100111000;
				8'b1000110: c <= 9'b100010111;
				8'b1110010: c <= 9'b1010101;
				8'b1010000: c <= 9'b101010010;
				8'b1111010: c <= 9'b100000100;
				8'b1010101: c <= 9'b110010011;
				8'b111011: c <= 9'b100101101;
				8'b1001101: c <= 9'b101001000;
				8'b111111: c <= 9'b10101001;
				8'b1101110: c <= 9'b101101010;
				8'b1111011: c <= 9'b100010001;
				8'b1001011: c <= 9'b101010;
				8'b1101111: c <= 9'b100001;
				8'b1101000: c <= 9'b100101000;
				8'b101100: c <= 9'b110001101;
				8'b100100: c <= 9'b111001110;
				8'b1111000: c <= 9'b111111101;
				8'b1000101: c <= 9'b100101010;
				8'b1011001: c <= 9'b10110011;
				8'b110100: c <= 9'b100100000;
				8'b1111001: c <= 9'b101010110;
				8'b1110001: c <= 9'b110110110;
				8'b1001111: c <= 9'b11001100;
				8'b1100101: c <= 9'b11001010;
				8'b1111110: c <= 9'b111101110;
				8'b1111100: c <= 9'b101010011;
				8'b1010110: c <= 9'b101101011;
				8'b110010: c <= 9'b11000001;
				8'b1101101: c <= 9'b111101110;
				8'b100011: c <= 9'b110110010;
				8'b1110101: c <= 9'b100010011;
				8'b1111101: c <= 9'b100111101;
				8'b101001: c <= 9'b100010;
				8'b1010010: c <= 9'b1001001;
				8'b1011000: c <= 9'b1110000;
				8'b101110: c <= 9'b100111010;
				8'b1000001: c <= 9'b110011100;
				default: c <= 9'b0;
			endcase
			9'b111000101 : case(di)
				8'b1000011: c <= 9'b111110011;
				8'b101000: c <= 9'b111011101;
				8'b111010: c <= 9'b10000111;
				8'b110110: c <= 9'b100101011;
				8'b1100100: c <= 9'b111101101;
				8'b1000000: c <= 9'b111101100;
				8'b1110110: c <= 9'b100011001;
				8'b100101: c <= 9'b10001010;
				8'b101111: c <= 9'b100110;
				8'b100110: c <= 9'b110000;
				8'b1100011: c <= 9'b111100010;
				8'b1001000: c <= 9'b101110001;
				8'b111000: c <= 9'b10010011;
				8'b110001: c <= 9'b100010001;
				8'b1010111: c <= 9'b100111010;
				8'b1001110: c <= 9'b101110;
				8'b1101010: c <= 9'b10111101;
				8'b1001001: c <= 9'b101111110;
				8'b1100000: c <= 9'b100001100;
				8'b110111: c <= 9'b11111010;
				8'b1011101: c <= 9'b11000001;
				8'b1011011: c <= 9'b11100011;
				8'b111001: c <= 9'b101011101;
				8'b1001010: c <= 9'b10010;
				8'b110011: c <= 9'b10010100;
				8'b1101100: c <= 9'b11110101;
				8'b1110111: c <= 9'b100001111;
				8'b101011: c <= 9'b1100001;
				8'b1101011: c <= 9'b111111101;
				8'b111100: c <= 9'b110110110;
				8'b1000111: c <= 9'b1111011;
				8'b1011111: c <= 9'b101101100;
				8'b1110100: c <= 9'b1000110;
				8'b101101: c <= 9'b110001101;
				8'b1010011: c <= 9'b100010110;
				8'b1100001: c <= 9'b110111010;
				8'b110101: c <= 9'b10111100;
				8'b1000100: c <= 9'b111001101;
				8'b1010001: c <= 9'b101111001;
				8'b1010100: c <= 9'b10001001;
				8'b1100110: c <= 9'b111111010;
				8'b101010: c <= 9'b10011010;
				8'b1011110: c <= 9'b100110100;
				8'b1100111: c <= 9'b100001101;
				8'b1011010: c <= 9'b10110110;
				8'b1000010: c <= 9'b100010011;
				8'b111101: c <= 9'b11;
				8'b110000: c <= 9'b100011111;
				8'b111110: c <= 9'b101110011;
				8'b1100010: c <= 9'b11000111;
				8'b1110000: c <= 9'b100111101;
				8'b1101001: c <= 9'b11100110;
				8'b1110011: c <= 9'b1000;
				8'b1001100: c <= 9'b101000100;
				8'b100001: c <= 9'b111111110;
				8'b1000110: c <= 9'b100001011;
				8'b1110010: c <= 9'b11010000;
				8'b1010000: c <= 9'b1101001;
				8'b1111010: c <= 9'b110111111;
				8'b1010101: c <= 9'b10000000;
				8'b111011: c <= 9'b100111110;
				8'b1001101: c <= 9'b101001000;
				8'b111111: c <= 9'b11010000;
				8'b1101110: c <= 9'b100110011;
				8'b1111011: c <= 9'b10011111;
				8'b1001011: c <= 9'b10100000;
				8'b1101111: c <= 9'b100001010;
				8'b1101000: c <= 9'b111101001;
				8'b101100: c <= 9'b110101110;
				8'b100100: c <= 9'b100010110;
				8'b1111000: c <= 9'b100011100;
				8'b1000101: c <= 9'b10110111;
				8'b1011001: c <= 9'b101000011;
				8'b110100: c <= 9'b100000001;
				8'b1111001: c <= 9'b110001000;
				8'b1110001: c <= 9'b110111010;
				8'b1001111: c <= 9'b11101;
				8'b1100101: c <= 9'b1111011;
				8'b1111110: c <= 9'b1000000;
				8'b1111100: c <= 9'b100100110;
				8'b1010110: c <= 9'b1111101;
				8'b110010: c <= 9'b10010011;
				8'b1101101: c <= 9'b100111011;
				8'b100011: c <= 9'b100101000;
				8'b1110101: c <= 9'b111000100;
				8'b1111101: c <= 9'b111111111;
				8'b101001: c <= 9'b100011100;
				8'b1010010: c <= 9'b101011001;
				8'b1011000: c <= 9'b100011010;
				8'b101110: c <= 9'b11001000;
				8'b1000001: c <= 9'b100010100;
				default: c <= 9'b0;
			endcase
			9'b110011000 : case(di)
				8'b1000011: c <= 9'b100011100;
				8'b101000: c <= 9'b110000;
				8'b111010: c <= 9'b1100110;
				8'b110110: c <= 9'b110001110;
				8'b1100100: c <= 9'b11011110;
				8'b1000000: c <= 9'b1001001;
				8'b1110110: c <= 9'b1100111;
				8'b100101: c <= 9'b10111000;
				8'b101111: c <= 9'b111000111;
				8'b100110: c <= 9'b100110110;
				8'b1100011: c <= 9'b110110110;
				8'b1001000: c <= 9'b11011110;
				8'b111000: c <= 9'b101011000;
				8'b110001: c <= 9'b11001011;
				8'b1010111: c <= 9'b111010110;
				8'b1001110: c <= 9'b110110000;
				8'b1101010: c <= 9'b111000100;
				8'b1001001: c <= 9'b110110100;
				8'b1100000: c <= 9'b101110110;
				8'b110111: c <= 9'b11010111;
				8'b1011101: c <= 9'b10001110;
				8'b1011011: c <= 9'b110101101;
				8'b111001: c <= 9'b110111001;
				8'b1001010: c <= 9'b110001000;
				8'b110011: c <= 9'b111001011;
				8'b1101100: c <= 9'b111000010;
				8'b1110111: c <= 9'b11010;
				8'b101011: c <= 9'b1101101;
				8'b1101011: c <= 9'b101001;
				8'b111100: c <= 9'b110101100;
				8'b1000111: c <= 9'b100110010;
				8'b1011111: c <= 9'b10101;
				8'b1110100: c <= 9'b100100011;
				8'b101101: c <= 9'b10011111;
				8'b1010011: c <= 9'b110110;
				8'b1100001: c <= 9'b101110;
				8'b110101: c <= 9'b10111110;
				8'b1000100: c <= 9'b111011011;
				8'b1010001: c <= 9'b10111000;
				8'b1010100: c <= 9'b100011111;
				8'b1100110: c <= 9'b11101;
				8'b101010: c <= 9'b111100001;
				8'b1011110: c <= 9'b110111000;
				8'b1100111: c <= 9'b111001011;
				8'b1011010: c <= 9'b10111110;
				8'b1000010: c <= 9'b101100011;
				8'b111101: c <= 9'b100011111;
				8'b110000: c <= 9'b101001100;
				8'b111110: c <= 9'b111011011;
				8'b1100010: c <= 9'b11001010;
				8'b1110000: c <= 9'b100100000;
				8'b1101001: c <= 9'b110010110;
				8'b1110011: c <= 9'b110001011;
				8'b1001100: c <= 9'b1011111;
				8'b100001: c <= 9'b111001110;
				8'b1000110: c <= 9'b1111011;
				8'b1110010: c <= 9'b1000010;
				8'b1010000: c <= 9'b111111101;
				8'b1111010: c <= 9'b101110111;
				8'b1010101: c <= 9'b110110101;
				8'b111011: c <= 9'b110000010;
				8'b1001101: c <= 9'b11111001;
				8'b111111: c <= 9'b1000101;
				8'b1101110: c <= 9'b110100100;
				8'b1111011: c <= 9'b100000111;
				8'b1001011: c <= 9'b110110111;
				8'b1101111: c <= 9'b100101111;
				8'b1101000: c <= 9'b110011100;
				8'b101100: c <= 9'b101011010;
				8'b100100: c <= 9'b111001110;
				8'b1111000: c <= 9'b11001000;
				8'b1000101: c <= 9'b11001001;
				8'b1011001: c <= 9'b110110101;
				8'b110100: c <= 9'b100011010;
				8'b1111001: c <= 9'b10001100;
				8'b1110001: c <= 9'b101101110;
				8'b1001111: c <= 9'b10111110;
				8'b1100101: c <= 9'b100101000;
				8'b1111110: c <= 9'b101101;
				8'b1111100: c <= 9'b100100101;
				8'b1010110: c <= 9'b1101101;
				8'b110010: c <= 9'b110011010;
				8'b1101101: c <= 9'b11010100;
				8'b100011: c <= 9'b110101;
				8'b1110101: c <= 9'b1;
				8'b1111101: c <= 9'b1011100;
				8'b101001: c <= 9'b111111111;
				8'b1010010: c <= 9'b11011000;
				8'b1011000: c <= 9'b10010011;
				8'b101110: c <= 9'b1111111;
				8'b1000001: c <= 9'b1100001;
				default: c <= 9'b0;
			endcase
			9'b11101 : case(di)
				8'b1000011: c <= 9'b11011010;
				8'b101000: c <= 9'b101101100;
				8'b111010: c <= 9'b100111100;
				8'b110110: c <= 9'b10101100;
				8'b1100100: c <= 9'b10110100;
				8'b1000000: c <= 9'b101111001;
				8'b1110110: c <= 9'b1000;
				8'b100101: c <= 9'b100000100;
				8'b101111: c <= 9'b110110101;
				8'b100110: c <= 9'b1010110;
				8'b1100011: c <= 9'b110011101;
				8'b1001000: c <= 9'b10000110;
				8'b111000: c <= 9'b101010001;
				8'b110001: c <= 9'b110011101;
				8'b1010111: c <= 9'b111011011;
				8'b1001110: c <= 9'b111000101;
				8'b1101010: c <= 9'b10001000;
				8'b1001001: c <= 9'b100101011;
				8'b1100000: c <= 9'b11011100;
				8'b110111: c <= 9'b1001100;
				8'b1011101: c <= 9'b11000001;
				8'b1011011: c <= 9'b110000;
				8'b111001: c <= 9'b110010001;
				8'b1001010: c <= 9'b100010000;
				8'b110011: c <= 9'b1011100;
				8'b1101100: c <= 9'b11111101;
				8'b1110111: c <= 9'b11001011;
				8'b101011: c <= 9'b110110;
				8'b1101011: c <= 9'b1110010;
				8'b111100: c <= 9'b101000101;
				8'b1000111: c <= 9'b100000000;
				8'b1011111: c <= 9'b100110101;
				8'b1110100: c <= 9'b1000111;
				8'b101101: c <= 9'b10110110;
				8'b1010011: c <= 9'b11001111;
				8'b1100001: c <= 9'b1001100;
				8'b110101: c <= 9'b1111111;
				8'b1000100: c <= 9'b111101010;
				8'b1010001: c <= 9'b10111100;
				8'b1010100: c <= 9'b110111110;
				8'b1100110: c <= 9'b100100001;
				8'b101010: c <= 9'b100011000;
				8'b1011110: c <= 9'b10110101;
				8'b1100111: c <= 9'b110101001;
				8'b1011010: c <= 9'b111111;
				8'b1000010: c <= 9'b10000010;
				8'b111101: c <= 9'b101011111;
				8'b110000: c <= 9'b110001101;
				8'b111110: c <= 9'b11110111;
				8'b1100010: c <= 9'b111100;
				8'b1110000: c <= 9'b10101011;
				8'b1101001: c <= 9'b10000111;
				8'b1110011: c <= 9'b111010;
				8'b1001100: c <= 9'b11001011;
				8'b100001: c <= 9'b110100100;
				8'b1000110: c <= 9'b101101000;
				8'b1110010: c <= 9'b10001011;
				8'b1010000: c <= 9'b110001011;
				8'b1111010: c <= 9'b10001100;
				8'b1010101: c <= 9'b11100110;
				8'b111011: c <= 9'b110110000;
				8'b1001101: c <= 9'b110011000;
				8'b111111: c <= 9'b111100110;
				8'b1101110: c <= 9'b110110011;
				8'b1111011: c <= 9'b101110011;
				8'b1001011: c <= 9'b100000011;
				8'b1101111: c <= 9'b100100010;
				8'b1101000: c <= 9'b111111000;
				8'b101100: c <= 9'b110100110;
				8'b100100: c <= 9'b11110100;
				8'b1111000: c <= 9'b1010010;
				8'b1000101: c <= 9'b11011110;
				8'b1011001: c <= 9'b10110100;
				8'b110100: c <= 9'b10010;
				8'b1111001: c <= 9'b110011001;
				8'b1110001: c <= 9'b111011111;
				8'b1001111: c <= 9'b1101010;
				8'b1100101: c <= 9'b101;
				8'b1111110: c <= 9'b100101;
				8'b1111100: c <= 9'b110011001;
				8'b1010110: c <= 9'b1111111;
				8'b110010: c <= 9'b1100000;
				8'b1101101: c <= 9'b11000010;
				8'b100011: c <= 9'b110100001;
				8'b1110101: c <= 9'b1001;
				8'b1111101: c <= 9'b111110000;
				8'b101001: c <= 9'b100111001;
				8'b1010010: c <= 9'b110000000;
				8'b1011000: c <= 9'b111111101;
				8'b101110: c <= 9'b101111110;
				8'b1000001: c <= 9'b110000111;
				default: c <= 9'b0;
			endcase
			9'b111011010 : case(di)
				8'b1000011: c <= 9'b11101001;
				8'b101000: c <= 9'b1000;
				8'b111010: c <= 9'b11100110;
				8'b110110: c <= 9'b110100000;
				8'b1100100: c <= 9'b110100110;
				8'b1000000: c <= 9'b11100010;
				8'b1110110: c <= 9'b100010100;
				8'b100101: c <= 9'b111000111;
				8'b101111: c <= 9'b111101;
				8'b100110: c <= 9'b10000011;
				8'b1100011: c <= 9'b100100000;
				8'b1001000: c <= 9'b1100010;
				8'b111000: c <= 9'b110000111;
				8'b110001: c <= 9'b101101000;
				8'b1010111: c <= 9'b100111100;
				8'b1001110: c <= 9'b111010010;
				8'b1101010: c <= 9'b110100011;
				8'b1001001: c <= 9'b111000000;
				8'b1100000: c <= 9'b10;
				8'b110111: c <= 9'b110100101;
				8'b1011101: c <= 9'b11010100;
				8'b1011011: c <= 9'b10111111;
				8'b111001: c <= 9'b11110110;
				8'b1001010: c <= 9'b100101000;
				8'b110011: c <= 9'b101100011;
				8'b1101100: c <= 9'b111100010;
				8'b1110111: c <= 9'b101011;
				8'b101011: c <= 9'b11111011;
				8'b1101011: c <= 9'b11001000;
				8'b111100: c <= 9'b111101101;
				8'b1000111: c <= 9'b110111011;
				8'b1011111: c <= 9'b11111;
				8'b1110100: c <= 9'b111100010;
				8'b101101: c <= 9'b101100101;
				8'b1010011: c <= 9'b1000;
				8'b1100001: c <= 9'b110100011;
				8'b110101: c <= 9'b110011010;
				8'b1000100: c <= 9'b110;
				8'b1010001: c <= 9'b101001111;
				8'b1010100: c <= 9'b111000110;
				8'b1100110: c <= 9'b100101101;
				8'b101010: c <= 9'b100110000;
				8'b1011110: c <= 9'b111010111;
				8'b1100111: c <= 9'b110001110;
				8'b1011010: c <= 9'b100011100;
				8'b1000010: c <= 9'b11100000;
				8'b111101: c <= 9'b11000000;
				8'b110000: c <= 9'b10101;
				8'b111110: c <= 9'b111001;
				8'b1100010: c <= 9'b100010010;
				8'b1110000: c <= 9'b100101;
				8'b1101001: c <= 9'b101101000;
				8'b1110011: c <= 9'b110111011;
				8'b1001100: c <= 9'b100011100;
				8'b100001: c <= 9'b11100000;
				8'b1000110: c <= 9'b1101000;
				8'b1110010: c <= 9'b111100;
				8'b1010000: c <= 9'b100000111;
				8'b1111010: c <= 9'b100111000;
				8'b1010101: c <= 9'b10001011;
				8'b111011: c <= 9'b110000011;
				8'b1001101: c <= 9'b11100001;
				8'b111111: c <= 9'b1111011;
				8'b1101110: c <= 9'b11101101;
				8'b1111011: c <= 9'b1110100;
				8'b1001011: c <= 9'b101000010;
				8'b1101111: c <= 9'b1011111;
				8'b1101000: c <= 9'b100110110;
				8'b101100: c <= 9'b1110001;
				8'b100100: c <= 9'b110010111;
				8'b1111000: c <= 9'b1101010;
				8'b1000101: c <= 9'b10101000;
				8'b1011001: c <= 9'b100000100;
				8'b110100: c <= 9'b11000;
				8'b1111001: c <= 9'b1101001;
				8'b1110001: c <= 9'b11110011;
				8'b1001111: c <= 9'b110101;
				8'b1100101: c <= 9'b10110;
				8'b1111110: c <= 9'b1010010;
				8'b1111100: c <= 9'b10110;
				8'b1010110: c <= 9'b100010111;
				8'b110010: c <= 9'b11011101;
				8'b1101101: c <= 9'b111100110;
				8'b100011: c <= 9'b111111111;
				8'b1110101: c <= 9'b111110011;
				8'b1111101: c <= 9'b110110111;
				8'b101001: c <= 9'b10110010;
				8'b1010010: c <= 9'b100100001;
				8'b1011000: c <= 9'b11100100;
				8'b101110: c <= 9'b1001;
				8'b1000001: c <= 9'b10000000;
				default: c <= 9'b0;
			endcase
			9'b101110011 : case(di)
				8'b1000011: c <= 9'b110010011;
				8'b101000: c <= 9'b11101011;
				8'b111010: c <= 9'b1001110;
				8'b110110: c <= 9'b101011001;
				8'b1100100: c <= 9'b110000;
				8'b1000000: c <= 9'b111000101;
				8'b1110110: c <= 9'b111011;
				8'b100101: c <= 9'b110011;
				8'b101111: c <= 9'b10000110;
				8'b100110: c <= 9'b100101001;
				8'b1100011: c <= 9'b111010100;
				8'b1001000: c <= 9'b110101010;
				8'b111000: c <= 9'b101111010;
				8'b110001: c <= 9'b1;
				8'b1010111: c <= 9'b111110011;
				8'b1001110: c <= 9'b101100111;
				8'b1101010: c <= 9'b10010101;
				8'b1001001: c <= 9'b10111110;
				8'b1100000: c <= 9'b1000110;
				8'b110111: c <= 9'b111101110;
				8'b1011101: c <= 9'b111010;
				8'b1011011: c <= 9'b110111;
				8'b111001: c <= 9'b10110111;
				8'b1001010: c <= 9'b100010000;
				8'b110011: c <= 9'b100110111;
				8'b1101100: c <= 9'b10101011;
				8'b1110111: c <= 9'b100010101;
				8'b101011: c <= 9'b101011101;
				8'b1101011: c <= 9'b110001101;
				8'b111100: c <= 9'b100000100;
				8'b1000111: c <= 9'b10010001;
				8'b1011111: c <= 9'b101100000;
				8'b1110100: c <= 9'b110111110;
				8'b101101: c <= 9'b10101001;
				8'b1010011: c <= 9'b10111010;
				8'b1100001: c <= 9'b100001001;
				8'b110101: c <= 9'b100;
				8'b1000100: c <= 9'b11000000;
				8'b1010001: c <= 9'b1110100;
				8'b1010100: c <= 9'b111110001;
				8'b1100110: c <= 9'b111011101;
				8'b101010: c <= 9'b111110101;
				8'b1011110: c <= 9'b101000111;
				8'b1100111: c <= 9'b101000011;
				8'b1011010: c <= 9'b11111101;
				8'b1000010: c <= 9'b10110001;
				8'b111101: c <= 9'b100000111;
				8'b110000: c <= 9'b1011001;
				8'b111110: c <= 9'b10011000;
				8'b1100010: c <= 9'b111111000;
				8'b1110000: c <= 9'b10011010;
				8'b1101001: c <= 9'b100101111;
				8'b1110011: c <= 9'b110;
				8'b1001100: c <= 9'b110111110;
				8'b100001: c <= 9'b100011100;
				8'b1000110: c <= 9'b111001100;
				8'b1110010: c <= 9'b110110101;
				8'b1010000: c <= 9'b100110011;
				8'b1111010: c <= 9'b10110110;
				8'b1010101: c <= 9'b11010111;
				8'b111011: c <= 9'b1111001;
				8'b1001101: c <= 9'b1100001;
				8'b111111: c <= 9'b10001110;
				8'b1101110: c <= 9'b10101011;
				8'b1111011: c <= 9'b111111101;
				8'b1001011: c <= 9'b11101;
				8'b1101111: c <= 9'b111110110;
				8'b1101000: c <= 9'b1000000;
				8'b101100: c <= 9'b111000010;
				8'b100100: c <= 9'b110100000;
				8'b1111000: c <= 9'b111000110;
				8'b1000101: c <= 9'b101000011;
				8'b1011001: c <= 9'b11111110;
				8'b110100: c <= 9'b11111011;
				8'b1111001: c <= 9'b10110101;
				8'b1110001: c <= 9'b100001100;
				8'b1001111: c <= 9'b1011010;
				8'b1100101: c <= 9'b100011100;
				8'b1111110: c <= 9'b10011000;
				8'b1111100: c <= 9'b101110111;
				8'b1010110: c <= 9'b10110110;
				8'b110010: c <= 9'b101001001;
				8'b1101101: c <= 9'b1101101;
				8'b100011: c <= 9'b1000111;
				8'b1110101: c <= 9'b110100000;
				8'b1111101: c <= 9'b11110100;
				8'b101001: c <= 9'b111001011;
				8'b1010010: c <= 9'b11001110;
				8'b1011000: c <= 9'b1010111;
				8'b101110: c <= 9'b11100101;
				8'b1000001: c <= 9'b11110100;
				default: c <= 9'b0;
			endcase
			9'b100000011 : case(di)
				8'b1000011: c <= 9'b111110101;
				8'b101000: c <= 9'b100101001;
				8'b111010: c <= 9'b1000011;
				8'b110110: c <= 9'b100010;
				8'b1100100: c <= 9'b111101000;
				8'b1000000: c <= 9'b101100111;
				8'b1110110: c <= 9'b10110001;
				8'b100101: c <= 9'b100001111;
				8'b101111: c <= 9'b100101111;
				8'b100110: c <= 9'b11101111;
				8'b1100011: c <= 9'b10001010;
				8'b1001000: c <= 9'b10010001;
				8'b111000: c <= 9'b111000010;
				8'b110001: c <= 9'b110101011;
				8'b1010111: c <= 9'b10011;
				8'b1001110: c <= 9'b11011010;
				8'b1101010: c <= 9'b10001001;
				8'b1001001: c <= 9'b111001010;
				8'b1100000: c <= 9'b100111101;
				8'b110111: c <= 9'b101001011;
				8'b1011101: c <= 9'b1001010;
				8'b1011011: c <= 9'b111011001;
				8'b111001: c <= 9'b10101101;
				8'b1001010: c <= 9'b1001001;
				8'b110011: c <= 9'b101011000;
				8'b1101100: c <= 9'b10111000;
				8'b1110111: c <= 9'b111110000;
				8'b101011: c <= 9'b1100011;
				8'b1101011: c <= 9'b101100011;
				8'b111100: c <= 9'b10111011;
				8'b1000111: c <= 9'b10000111;
				8'b1011111: c <= 9'b101010000;
				8'b1110100: c <= 9'b11001110;
				8'b101101: c <= 9'b100101100;
				8'b1010011: c <= 9'b110011000;
				8'b1100001: c <= 9'b101101111;
				8'b110101: c <= 9'b110001110;
				8'b1000100: c <= 9'b100100010;
				8'b1010001: c <= 9'b101110000;
				8'b1010100: c <= 9'b101100010;
				8'b1100110: c <= 9'b11011110;
				8'b101010: c <= 9'b10001001;
				8'b1011110: c <= 9'b110101100;
				8'b1100111: c <= 9'b101100100;
				8'b1011010: c <= 9'b100100110;
				8'b1000010: c <= 9'b100010010;
				8'b111101: c <= 9'b10100101;
				8'b110000: c <= 9'b111111010;
				8'b111110: c <= 9'b1101010;
				8'b1100010: c <= 9'b10101111;
				8'b1110000: c <= 9'b111001111;
				8'b1101001: c <= 9'b1111110;
				8'b1110011: c <= 9'b101111111;
				8'b1001100: c <= 9'b110101001;
				8'b100001: c <= 9'b110100110;
				8'b1000110: c <= 9'b101110110;
				8'b1110010: c <= 9'b1010011;
				8'b1010000: c <= 9'b101;
				8'b1111010: c <= 9'b111100011;
				8'b1010101: c <= 9'b101011111;
				8'b111011: c <= 9'b11010001;
				8'b1001101: c <= 9'b100010001;
				8'b111111: c <= 9'b11100;
				8'b1101110: c <= 9'b1110100;
				8'b1111011: c <= 9'b11111010;
				8'b1001011: c <= 9'b10101011;
				8'b1101111: c <= 9'b100010;
				8'b1101000: c <= 9'b10011000;
				8'b101100: c <= 9'b1011011;
				8'b100100: c <= 9'b110011100;
				8'b1111000: c <= 9'b11010000;
				8'b1000101: c <= 9'b111001010;
				8'b1011001: c <= 9'b100111001;
				8'b110100: c <= 9'b100001011;
				8'b1111001: c <= 9'b110001011;
				8'b1110001: c <= 9'b111101000;
				8'b1001111: c <= 9'b11111011;
				8'b1100101: c <= 9'b110001100;
				8'b1111110: c <= 9'b100000011;
				8'b1111100: c <= 9'b100111011;
				8'b1010110: c <= 9'b101000010;
				8'b110010: c <= 9'b1001001;
				8'b1101101: c <= 9'b10011011;
				8'b100011: c <= 9'b111011010;
				8'b1110101: c <= 9'b10000000;
				8'b1111101: c <= 9'b110100;
				8'b101001: c <= 9'b1111110;
				8'b1010010: c <= 9'b100000001;
				8'b1011000: c <= 9'b10101010;
				8'b101110: c <= 9'b100110110;
				8'b1000001: c <= 9'b100010101;
				default: c <= 9'b0;
			endcase
			9'b1001001 : case(di)
				8'b1000011: c <= 9'b101001001;
				8'b101000: c <= 9'b11101001;
				8'b111010: c <= 9'b100000001;
				8'b110110: c <= 9'b1011100;
				8'b1100100: c <= 9'b1100000;
				8'b1000000: c <= 9'b10111101;
				8'b1110110: c <= 9'b110001010;
				8'b100101: c <= 9'b101100110;
				8'b101111: c <= 9'b101111111;
				8'b100110: c <= 9'b10001000;
				8'b1100011: c <= 9'b1011011;
				8'b1001000: c <= 9'b100101100;
				8'b111000: c <= 9'b11111011;
				8'b110001: c <= 9'b100001100;
				8'b1010111: c <= 9'b110110100;
				8'b1001110: c <= 9'b11001010;
				8'b1101010: c <= 9'b11101101;
				8'b1001001: c <= 9'b100001101;
				8'b1100000: c <= 9'b10001000;
				8'b110111: c <= 9'b110111010;
				8'b1011101: c <= 9'b10000000;
				8'b1011011: c <= 9'b100;
				8'b111001: c <= 9'b1011011;
				8'b1001010: c <= 9'b101011101;
				8'b110011: c <= 9'b110110100;
				8'b1101100: c <= 9'b10110011;
				8'b1110111: c <= 9'b1111011;
				8'b101011: c <= 9'b111010;
				8'b1101011: c <= 9'b100001111;
				8'b111100: c <= 9'b1110100;
				8'b1000111: c <= 9'b11000000;
				8'b1011111: c <= 9'b100011;
				8'b1110100: c <= 9'b10101100;
				8'b101101: c <= 9'b1110111;
				8'b1010011: c <= 9'b100110;
				8'b1100001: c <= 9'b110010100;
				8'b110101: c <= 9'b10011011;
				8'b1000100: c <= 9'b111101000;
				8'b1010001: c <= 9'b1000011;
				8'b1010100: c <= 9'b110100110;
				8'b1100110: c <= 9'b1101101;
				8'b101010: c <= 9'b100101110;
				8'b1011110: c <= 9'b101111111;
				8'b1100111: c <= 9'b100101011;
				8'b1011010: c <= 9'b110100111;
				8'b1000010: c <= 9'b1100;
				8'b111101: c <= 9'b1111;
				8'b110000: c <= 9'b1111111;
				8'b111110: c <= 9'b1011011;
				8'b1100010: c <= 9'b1101100;
				8'b1110000: c <= 9'b10011010;
				8'b1101001: c <= 9'b10010;
				8'b1110011: c <= 9'b11001;
				8'b1001100: c <= 9'b110101;
				8'b100001: c <= 9'b10011011;
				8'b1000110: c <= 9'b100100011;
				8'b1110010: c <= 9'b1010001;
				8'b1010000: c <= 9'b101001111;
				8'b1111010: c <= 9'b100011010;
				8'b1010101: c <= 9'b100011000;
				8'b111011: c <= 9'b111000011;
				8'b1001101: c <= 9'b11111000;
				8'b111111: c <= 9'b11110000;
				8'b1101110: c <= 9'b100000000;
				8'b1111011: c <= 9'b10100;
				8'b1001011: c <= 9'b11001110;
				8'b1101111: c <= 9'b101;
				8'b1101000: c <= 9'b101010000;
				8'b101100: c <= 9'b11101;
				8'b100100: c <= 9'b11101011;
				8'b1111000: c <= 9'b100111100;
				8'b1000101: c <= 9'b11000000;
				8'b1011001: c <= 9'b1111101;
				8'b110100: c <= 9'b1001110;
				8'b1111001: c <= 9'b101110110;
				8'b1110001: c <= 9'b110100101;
				8'b1001111: c <= 9'b111111;
				8'b1100101: c <= 9'b10110011;
				8'b1111110: c <= 9'b111011100;
				8'b1111100: c <= 9'b101110010;
				8'b1010110: c <= 9'b10010110;
				8'b110010: c <= 9'b110011110;
				8'b1101101: c <= 9'b101101111;
				8'b100011: c <= 9'b111100110;
				8'b1110101: c <= 9'b100101000;
				8'b1111101: c <= 9'b101101;
				8'b101001: c <= 9'b111011111;
				8'b1010010: c <= 9'b1110000;
				8'b1011000: c <= 9'b100101111;
				8'b101110: c <= 9'b110011011;
				8'b1000001: c <= 9'b111000010;
				default: c <= 9'b0;
			endcase
			9'b1101100 : case(di)
				8'b1000011: c <= 9'b101000;
				8'b101000: c <= 9'b101000111;
				8'b111010: c <= 9'b10101011;
				8'b110110: c <= 9'b11001111;
				8'b1100100: c <= 9'b111110000;
				8'b1000000: c <= 9'b110001100;
				8'b1110110: c <= 9'b100101100;
				8'b100101: c <= 9'b111010000;
				8'b101111: c <= 9'b100000010;
				8'b100110: c <= 9'b10111;
				8'b1100011: c <= 9'b10011;
				8'b1001000: c <= 9'b10111110;
				8'b111000: c <= 9'b110000;
				8'b110001: c <= 9'b110000101;
				8'b1010111: c <= 9'b10000111;
				8'b1001110: c <= 9'b101100111;
				8'b1101010: c <= 9'b11010011;
				8'b1001001: c <= 9'b110011011;
				8'b1100000: c <= 9'b101101011;
				8'b110111: c <= 9'b11001101;
				8'b1011101: c <= 9'b1011010;
				8'b1011011: c <= 9'b101110100;
				8'b111001: c <= 9'b101111000;
				8'b1001010: c <= 9'b101010010;
				8'b110011: c <= 9'b1101110;
				8'b1101100: c <= 9'b111011010;
				8'b1110111: c <= 9'b100101111;
				8'b101011: c <= 9'b101001;
				8'b1101011: c <= 9'b110111011;
				8'b111100: c <= 9'b1111010;
				8'b1000111: c <= 9'b110011110;
				8'b1011111: c <= 9'b111;
				8'b1110100: c <= 9'b10101;
				8'b101101: c <= 9'b111100110;
				8'b1010011: c <= 9'b110100011;
				8'b1100001: c <= 9'b100111101;
				8'b110101: c <= 9'b111011100;
				8'b1000100: c <= 9'b101110100;
				8'b1010001: c <= 9'b111100010;
				8'b1010100: c <= 9'b111111101;
				8'b1100110: c <= 9'b100101010;
				8'b101010: c <= 9'b101001111;
				8'b1011110: c <= 9'b100000100;
				8'b1100111: c <= 9'b11001101;
				8'b1011010: c <= 9'b1111010;
				8'b1000010: c <= 9'b11101;
				8'b111101: c <= 9'b110000110;
				8'b110000: c <= 9'b1111000;
				8'b111110: c <= 9'b100100110;
				8'b1100010: c <= 9'b101001111;
				8'b1110000: c <= 9'b1100011;
				8'b1101001: c <= 9'b10010001;
				8'b1110011: c <= 9'b100100011;
				8'b1001100: c <= 9'b11001001;
				8'b100001: c <= 9'b10110101;
				8'b1000110: c <= 9'b110111110;
				8'b1110010: c <= 9'b1000110;
				8'b1010000: c <= 9'b101110011;
				8'b1111010: c <= 9'b101011000;
				8'b1010101: c <= 9'b111000111;
				8'b111011: c <= 9'b101111111;
				8'b1001101: c <= 9'b111000000;
				8'b111111: c <= 9'b111;
				8'b1101110: c <= 9'b11001110;
				8'b1111011: c <= 9'b101100000;
				8'b1001011: c <= 9'b11010011;
				8'b1101111: c <= 9'b10000101;
				8'b1101000: c <= 9'b101101010;
				8'b101100: c <= 9'b100011011;
				8'b100100: c <= 9'b1000010;
				8'b1111000: c <= 9'b110010011;
				8'b1000101: c <= 9'b100110010;
				8'b1011001: c <= 9'b110101010;
				8'b110100: c <= 9'b1001011;
				8'b1111001: c <= 9'b101001;
				8'b1110001: c <= 9'b111111010;
				8'b1001111: c <= 9'b1101;
				8'b1100101: c <= 9'b10000110;
				8'b1111110: c <= 9'b11110001;
				8'b1111100: c <= 9'b111001;
				8'b1010110: c <= 9'b100111110;
				8'b110010: c <= 9'b10010101;
				8'b1101101: c <= 9'b110010;
				8'b100011: c <= 9'b111101101;
				8'b1110101: c <= 9'b11101111;
				8'b1111101: c <= 9'b10111001;
				8'b101001: c <= 9'b111000111;
				8'b1010010: c <= 9'b11111011;
				8'b1011000: c <= 9'b100010101;
				8'b101110: c <= 9'b101001001;
				8'b1000001: c <= 9'b110111010;
				default: c <= 9'b0;
			endcase
			9'b11101100 : case(di)
				8'b1000011: c <= 9'b1000110;
				8'b101000: c <= 9'b110110111;
				8'b111010: c <= 9'b101000001;
				8'b110110: c <= 9'b11110110;
				8'b1100100: c <= 9'b110101100;
				8'b1000000: c <= 9'b11000110;
				8'b1110110: c <= 9'b111010100;
				8'b100101: c <= 9'b111001111;
				8'b101111: c <= 9'b111111101;
				8'b100110: c <= 9'b111001011;
				8'b1100011: c <= 9'b110101101;
				8'b1001000: c <= 9'b111001010;
				8'b111000: c <= 9'b100101010;
				8'b110001: c <= 9'b111000010;
				8'b1010111: c <= 9'b110001010;
				8'b1001110: c <= 9'b10111;
				8'b1101010: c <= 9'b10111110;
				8'b1001001: c <= 9'b10000000;
				8'b1100000: c <= 9'b10100011;
				8'b110111: c <= 9'b100100;
				8'b1011101: c <= 9'b11110000;
				8'b1011011: c <= 9'b101010101;
				8'b111001: c <= 9'b110011110;
				8'b1001010: c <= 9'b1000101;
				8'b110011: c <= 9'b111000000;
				8'b1101100: c <= 9'b101110;
				8'b1110111: c <= 9'b110000;
				8'b101011: c <= 9'b11110110;
				8'b1101011: c <= 9'b11111011;
				8'b111100: c <= 9'b111100010;
				8'b1000111: c <= 9'b101100001;
				8'b1011111: c <= 9'b100010111;
				8'b1110100: c <= 9'b100000101;
				8'b101101: c <= 9'b110010100;
				8'b1010011: c <= 9'b100101010;
				8'b1100001: c <= 9'b100000000;
				8'b110101: c <= 9'b101100011;
				8'b1000100: c <= 9'b101011011;
				8'b1010001: c <= 9'b11001;
				8'b1010100: c <= 9'b11110100;
				8'b1100110: c <= 9'b1100110;
				8'b101010: c <= 9'b110110000;
				8'b1011110: c <= 9'b11100110;
				8'b1100111: c <= 9'b111001010;
				8'b1011010: c <= 9'b1000110;
				8'b1000010: c <= 9'b11100110;
				8'b111101: c <= 9'b100001101;
				8'b110000: c <= 9'b10110;
				8'b111110: c <= 9'b11011101;
				8'b1100010: c <= 9'b110100100;
				8'b1110000: c <= 9'b111;
				8'b1101001: c <= 9'b110000;
				8'b1110011: c <= 9'b100011101;
				8'b1001100: c <= 9'b101111111;
				8'b100001: c <= 9'b111110101;
				8'b1000110: c <= 9'b11111;
				8'b1110010: c <= 9'b111100111;
				8'b1010000: c <= 9'b101101000;
				8'b1111010: c <= 9'b1011011;
				8'b1010101: c <= 9'b100111;
				8'b111011: c <= 9'b100101100;
				8'b1001101: c <= 9'b101000010;
				8'b111111: c <= 9'b101000100;
				8'b1101110: c <= 9'b100101010;
				8'b1111011: c <= 9'b101011;
				8'b1001011: c <= 9'b100010111;
				8'b1101111: c <= 9'b10011001;
				8'b1101000: c <= 9'b11110;
				8'b101100: c <= 9'b110111010;
				8'b100100: c <= 9'b100010111;
				8'b1111000: c <= 9'b100000001;
				8'b1000101: c <= 9'b11110;
				8'b1011001: c <= 9'b101101110;
				8'b110100: c <= 9'b1000;
				8'b1111001: c <= 9'b1000101;
				8'b1110001: c <= 9'b10101011;
				8'b1001111: c <= 9'b111111;
				8'b1100101: c <= 9'b1000111;
				8'b1111110: c <= 9'b1011001;
				8'b1111100: c <= 9'b10000111;
				8'b1010110: c <= 9'b100011100;
				8'b110010: c <= 9'b10000000;
				8'b1101101: c <= 9'b11011010;
				8'b100011: c <= 9'b110000101;
				8'b1110101: c <= 9'b10001001;
				8'b1111101: c <= 9'b111001010;
				8'b101001: c <= 9'b1010111;
				8'b1010010: c <= 9'b111000010;
				8'b1011000: c <= 9'b100011011;
				8'b101110: c <= 9'b11111001;
				8'b1000001: c <= 9'b1100101;
				default: c <= 9'b0;
			endcase
			9'b101000101 : case(di)
				8'b1000011: c <= 9'b10001111;
				8'b101000: c <= 9'b111001000;
				8'b111010: c <= 9'b10001011;
				8'b110110: c <= 9'b100011011;
				8'b1100100: c <= 9'b100100111;
				8'b1000000: c <= 9'b10000011;
				8'b1110110: c <= 9'b100000011;
				8'b100101: c <= 9'b101001100;
				8'b101111: c <= 9'b101001;
				8'b100110: c <= 9'b110011001;
				8'b1100011: c <= 9'b1110010;
				8'b1001000: c <= 9'b11010111;
				8'b111000: c <= 9'b10101101;
				8'b110001: c <= 9'b1010011;
				8'b1010111: c <= 9'b1010001;
				8'b1001110: c <= 9'b10110010;
				8'b1101010: c <= 9'b10010011;
				8'b1001001: c <= 9'b1010001;
				8'b1100000: c <= 9'b1111110;
				8'b110111: c <= 9'b10000010;
				8'b1011101: c <= 9'b111101110;
				8'b1011011: c <= 9'b100010110;
				8'b111001: c <= 9'b110011001;
				8'b1001010: c <= 9'b11000010;
				8'b110011: c <= 9'b11010;
				8'b1101100: c <= 9'b11000100;
				8'b1110111: c <= 9'b111000;
				8'b101011: c <= 9'b100101110;
				8'b1101011: c <= 9'b111011110;
				8'b111100: c <= 9'b111011010;
				8'b1000111: c <= 9'b1101001;
				8'b1011111: c <= 9'b11110011;
				8'b1110100: c <= 9'b100010010;
				8'b101101: c <= 9'b1101110;
				8'b1010011: c <= 9'b110001010;
				8'b1100001: c <= 9'b11100011;
				8'b110101: c <= 9'b10011010;
				8'b1000100: c <= 9'b10010;
				8'b1010001: c <= 9'b110001111;
				8'b1010100: c <= 9'b11001001;
				8'b1100110: c <= 9'b1001010;
				8'b101010: c <= 9'b110010001;
				8'b1011110: c <= 9'b101100000;
				8'b1100111: c <= 9'b110;
				8'b1011010: c <= 9'b10100101;
				8'b1000010: c <= 9'b111001010;
				8'b111101: c <= 9'b111011111;
				8'b110000: c <= 9'b100111000;
				8'b111110: c <= 9'b101011110;
				8'b1100010: c <= 9'b110;
				8'b1110000: c <= 9'b11001000;
				8'b1101001: c <= 9'b1011010;
				8'b1110011: c <= 9'b110010001;
				8'b1001100: c <= 9'b110101100;
				8'b100001: c <= 9'b1100001;
				8'b1000110: c <= 9'b1101111;
				8'b1110010: c <= 9'b100000011;
				8'b1010000: c <= 9'b110001101;
				8'b1111010: c <= 9'b10110;
				8'b1010101: c <= 9'b11100111;
				8'b111011: c <= 9'b101110000;
				8'b1001101: c <= 9'b11001;
				8'b111111: c <= 9'b101001110;
				8'b1101110: c <= 9'b10001110;
				8'b1111011: c <= 9'b10000101;
				8'b1001011: c <= 9'b111000000;
				8'b1101111: c <= 9'b110110010;
				8'b1101000: c <= 9'b111000010;
				8'b101100: c <= 9'b10001001;
				8'b100100: c <= 9'b11000010;
				8'b1111000: c <= 9'b1110101;
				8'b1000101: c <= 9'b1100010;
				8'b1011001: c <= 9'b1101010;
				8'b110100: c <= 9'b110001110;
				8'b1111001: c <= 9'b111010001;
				8'b1110001: c <= 9'b1000100;
				8'b1001111: c <= 9'b101110101;
				8'b1100101: c <= 9'b10111011;
				8'b1111110: c <= 9'b101000010;
				8'b1111100: c <= 9'b100010010;
				8'b1010110: c <= 9'b11100;
				8'b110010: c <= 9'b100001;
				8'b1101101: c <= 9'b111000101;
				8'b100011: c <= 9'b101001010;
				8'b1110101: c <= 9'b11011110;
				8'b1111101: c <= 9'b110011001;
				8'b101001: c <= 9'b11000010;
				8'b1010010: c <= 9'b1110000;
				8'b1011000: c <= 9'b1101;
				8'b101110: c <= 9'b111101000;
				8'b1000001: c <= 9'b10100000;
				default: c <= 9'b0;
			endcase
			9'b110011101 : case(di)
				8'b1000011: c <= 9'b110100001;
				8'b101000: c <= 9'b110000;
				8'b111010: c <= 9'b111010110;
				8'b110110: c <= 9'b10001011;
				8'b1100100: c <= 9'b10000010;
				8'b1000000: c <= 9'b100000101;
				8'b1110110: c <= 9'b100011111;
				8'b100101: c <= 9'b100111011;
				8'b101111: c <= 9'b11010000;
				8'b100110: c <= 9'b1011;
				8'b1100011: c <= 9'b100000011;
				8'b1001000: c <= 9'b110000001;
				8'b111000: c <= 9'b101101010;
				8'b110001: c <= 9'b10101111;
				8'b1010111: c <= 9'b110010;
				8'b1001110: c <= 9'b11001100;
				8'b1101010: c <= 9'b1100000;
				8'b1001001: c <= 9'b111001010;
				8'b1100000: c <= 9'b101110010;
				8'b110111: c <= 9'b111111;
				8'b1011101: c <= 9'b11111011;
				8'b1011011: c <= 9'b1100010;
				8'b111001: c <= 9'b1011000;
				8'b1001010: c <= 9'b100010010;
				8'b110011: c <= 9'b100001011;
				8'b1101100: c <= 9'b1101000;
				8'b1110111: c <= 9'b10101111;
				8'b101011: c <= 9'b10001100;
				8'b1101011: c <= 9'b101000001;
				8'b111100: c <= 9'b110001101;
				8'b1000111: c <= 9'b101001111;
				8'b1011111: c <= 9'b10101111;
				8'b1110100: c <= 9'b1010010;
				8'b101101: c <= 9'b111100110;
				8'b1010011: c <= 9'b110110010;
				8'b1100001: c <= 9'b10100100;
				8'b110101: c <= 9'b10001000;
				8'b1000100: c <= 9'b101101000;
				8'b1010001: c <= 9'b11001010;
				8'b1010100: c <= 9'b110001000;
				8'b1100110: c <= 9'b110;
				8'b101010: c <= 9'b101010010;
				8'b1011110: c <= 9'b10000010;
				8'b1100111: c <= 9'b111101111;
				8'b1011010: c <= 9'b100111011;
				8'b1000010: c <= 9'b111111;
				8'b111101: c <= 9'b111000;
				8'b110000: c <= 9'b100000110;
				8'b111110: c <= 9'b100000011;
				8'b1100010: c <= 9'b110101100;
				8'b1110000: c <= 9'b10101011;
				8'b1101001: c <= 9'b111001011;
				8'b1110011: c <= 9'b111010100;
				8'b1001100: c <= 9'b100110101;
				8'b100001: c <= 9'b110110000;
				8'b1000110: c <= 9'b100010011;
				8'b1110010: c <= 9'b10001011;
				8'b1010000: c <= 9'b11100101;
				8'b1111010: c <= 9'b10111000;
				8'b1010101: c <= 9'b110000010;
				8'b111011: c <= 9'b111100100;
				8'b1001101: c <= 9'b1110000;
				8'b111111: c <= 9'b10101100;
				8'b1101110: c <= 9'b100100000;
				8'b1111011: c <= 9'b1000;
				8'b1001011: c <= 9'b100010000;
				8'b1101111: c <= 9'b110101100;
				8'b1101000: c <= 9'b11111100;
				8'b101100: c <= 9'b101110110;
				8'b100100: c <= 9'b111010000;
				8'b1111000: c <= 9'b11001001;
				8'b1000101: c <= 9'b110000111;
				8'b1011001: c <= 9'b111101000;
				8'b110100: c <= 9'b101110001;
				8'b1111001: c <= 9'b111011001;
				8'b1110001: c <= 9'b111100010;
				8'b1001111: c <= 9'b10010111;
				8'b1100101: c <= 9'b11000011;
				8'b1111110: c <= 9'b110000110;
				8'b1111100: c <= 9'b10011000;
				8'b1010110: c <= 9'b101101101;
				8'b110010: c <= 9'b101100101;
				8'b1101101: c <= 9'b10000110;
				8'b100011: c <= 9'b10100111;
				8'b1110101: c <= 9'b11101001;
				8'b1111101: c <= 9'b101;
				8'b101001: c <= 9'b100101011;
				8'b1010010: c <= 9'b10100010;
				8'b1011000: c <= 9'b100111111;
				8'b101110: c <= 9'b11001001;
				8'b1000001: c <= 9'b111011;
				default: c <= 9'b0;
			endcase
			9'b11101101 : case(di)
				8'b1000011: c <= 9'b110101001;
				8'b101000: c <= 9'b111010001;
				8'b111010: c <= 9'b11110;
				8'b110110: c <= 9'b100101000;
				8'b1100100: c <= 9'b111111110;
				8'b1000000: c <= 9'b100000111;
				8'b1110110: c <= 9'b100111110;
				8'b100101: c <= 9'b101101001;
				8'b101111: c <= 9'b101100100;
				8'b100110: c <= 9'b100000000;
				8'b1100011: c <= 9'b100111011;
				8'b1001000: c <= 9'b1101;
				8'b111000: c <= 9'b100000110;
				8'b110001: c <= 9'b10110001;
				8'b1010111: c <= 9'b11111010;
				8'b1001110: c <= 9'b110000101;
				8'b1101010: c <= 9'b110110000;
				8'b1001001: c <= 9'b10;
				8'b1100000: c <= 9'b101010111;
				8'b110111: c <= 9'b1111001;
				8'b1011101: c <= 9'b1010001;
				8'b1011011: c <= 9'b1101000;
				8'b111001: c <= 9'b110110010;
				8'b1001010: c <= 9'b11110001;
				8'b110011: c <= 9'b110100000;
				8'b1101100: c <= 9'b1110;
				8'b1110111: c <= 9'b111001010;
				8'b101011: c <= 9'b111011001;
				8'b1101011: c <= 9'b110111;
				8'b111100: c <= 9'b1000110;
				8'b1000111: c <= 9'b110100010;
				8'b1011111: c <= 9'b10001110;
				8'b1110100: c <= 9'b111111011;
				8'b101101: c <= 9'b101100010;
				8'b1010011: c <= 9'b10110011;
				8'b1100001: c <= 9'b111111110;
				8'b110101: c <= 9'b110001101;
				8'b1000100: c <= 9'b10011101;
				8'b1010001: c <= 9'b100000110;
				8'b1010100: c <= 9'b10010;
				8'b1100110: c <= 9'b1011010;
				8'b101010: c <= 9'b1000100;
				8'b1011110: c <= 9'b1010110;
				8'b1100111: c <= 9'b100101010;
				8'b1011010: c <= 9'b101101111;
				8'b1000010: c <= 9'b100001001;
				8'b111101: c <= 9'b11011100;
				8'b110000: c <= 9'b110000010;
				8'b111110: c <= 9'b111100100;
				8'b1100010: c <= 9'b110111001;
				8'b1110000: c <= 9'b10111100;
				8'b1101001: c <= 9'b111010;
				8'b1110011: c <= 9'b110000101;
				8'b1001100: c <= 9'b110011100;
				8'b100001: c <= 9'b100110101;
				8'b1000110: c <= 9'b11111110;
				8'b1110010: c <= 9'b1001010;
				8'b1010000: c <= 9'b100001110;
				8'b1111010: c <= 9'b10010111;
				8'b1010101: c <= 9'b111010000;
				8'b111011: c <= 9'b11101000;
				8'b1001101: c <= 9'b10000111;
				8'b111111: c <= 9'b101011001;
				8'b1101110: c <= 9'b110000101;
				8'b1111011: c <= 9'b110011111;
				8'b1001011: c <= 9'b101000101;
				8'b1101111: c <= 9'b101000111;
				8'b1101000: c <= 9'b1100100;
				8'b101100: c <= 9'b100001011;
				8'b100100: c <= 9'b101010111;
				8'b1111000: c <= 9'b101000110;
				8'b1000101: c <= 9'b110000;
				8'b1011001: c <= 9'b101111110;
				8'b110100: c <= 9'b110111110;
				8'b1111001: c <= 9'b1100;
				8'b1110001: c <= 9'b100011010;
				8'b1001111: c <= 9'b100111000;
				8'b1100101: c <= 9'b111001;
				8'b1111110: c <= 9'b1100010;
				8'b1111100: c <= 9'b111011010;
				8'b1010110: c <= 9'b111111010;
				8'b110010: c <= 9'b110000101;
				8'b1101101: c <= 9'b10010110;
				8'b100011: c <= 9'b110110101;
				8'b1110101: c <= 9'b110001100;
				8'b1111101: c <= 9'b10001111;
				8'b101001: c <= 9'b110100;
				8'b1010010: c <= 9'b10100111;
				8'b1011000: c <= 9'b11011110;
				8'b101110: c <= 9'b1011;
				8'b1000001: c <= 9'b101100;
				default: c <= 9'b0;
			endcase
			9'b101001001 : case(di)
				8'b1000011: c <= 9'b1110000;
				8'b101000: c <= 9'b10111101;
				8'b111010: c <= 9'b10100100;
				8'b110110: c <= 9'b111001001;
				8'b1100100: c <= 9'b100100101;
				8'b1000000: c <= 9'b110100100;
				8'b1110110: c <= 9'b10010110;
				8'b100101: c <= 9'b10010001;
				8'b101111: c <= 9'b111100110;
				8'b100110: c <= 9'b110110111;
				8'b1100011: c <= 9'b111111111;
				8'b1001000: c <= 9'b1011010;
				8'b111000: c <= 9'b100000010;
				8'b110001: c <= 9'b101000100;
				8'b1010111: c <= 9'b1100011;
				8'b1001110: c <= 9'b100100;
				8'b1101010: c <= 9'b101110100;
				8'b1001001: c <= 9'b101111110;
				8'b1100000: c <= 9'b11010;
				8'b110111: c <= 9'b100001010;
				8'b1011101: c <= 9'b1001110;
				8'b1011011: c <= 9'b110010101;
				8'b111001: c <= 9'b11110001;
				8'b1001010: c <= 9'b1111100;
				8'b110011: c <= 9'b101110001;
				8'b1101100: c <= 9'b11110000;
				8'b1110111: c <= 9'b100010010;
				8'b101011: c <= 9'b101101111;
				8'b1101011: c <= 9'b11011000;
				8'b111100: c <= 9'b11101;
				8'b1000111: c <= 9'b101110011;
				8'b1011111: c <= 9'b100010010;
				8'b1110100: c <= 9'b111001111;
				8'b101101: c <= 9'b100000010;
				8'b1010011: c <= 9'b100001100;
				8'b1100001: c <= 9'b110011101;
				8'b110101: c <= 9'b100111;
				8'b1000100: c <= 9'b111101001;
				8'b1010001: c <= 9'b110100111;
				8'b1010100: c <= 9'b11110110;
				8'b1100110: c <= 9'b110111110;
				8'b101010: c <= 9'b100011001;
				8'b1011110: c <= 9'b10110;
				8'b1100111: c <= 9'b1111011;
				8'b1011010: c <= 9'b1001110;
				8'b1000010: c <= 9'b100111;
				8'b111101: c <= 9'b10101101;
				8'b110000: c <= 9'b111111010;
				8'b111110: c <= 9'b110001000;
				8'b1100010: c <= 9'b11011110;
				8'b1110000: c <= 9'b1010000;
				8'b1101001: c <= 9'b110;
				8'b1110011: c <= 9'b101001011;
				8'b1001100: c <= 9'b100110101;
				8'b100001: c <= 9'b110011011;
				8'b1000110: c <= 9'b10001100;
				8'b1110010: c <= 9'b11110;
				8'b1010000: c <= 9'b11001100;
				8'b1111010: c <= 9'b100010000;
				8'b1010101: c <= 9'b111101110;
				8'b111011: c <= 9'b111011100;
				8'b1001101: c <= 9'b101100000;
				8'b111111: c <= 9'b1110;
				8'b1101110: c <= 9'b10001111;
				8'b1111011: c <= 9'b11;
				8'b1001011: c <= 9'b111011110;
				8'b1101111: c <= 9'b110100100;
				8'b1101000: c <= 9'b10011100;
				8'b101100: c <= 9'b1011011;
				8'b100100: c <= 9'b10101;
				8'b1111000: c <= 9'b101100000;
				8'b1000101: c <= 9'b1;
				8'b1011001: c <= 9'b101010001;
				8'b110100: c <= 9'b11110100;
				8'b1111001: c <= 9'b101010111;
				8'b1110001: c <= 9'b1011000;
				8'b1001111: c <= 9'b110001000;
				8'b1100101: c <= 9'b111110110;
				8'b1111110: c <= 9'b111100;
				8'b1111100: c <= 9'b110011;
				8'b1010110: c <= 9'b101000111;
				8'b110010: c <= 9'b100111101;
				8'b1101101: c <= 9'b100101010;
				8'b100011: c <= 9'b100110111;
				8'b1110101: c <= 9'b11110100;
				8'b1111101: c <= 9'b10010111;
				8'b101001: c <= 9'b100010101;
				8'b1010010: c <= 9'b10110111;
				8'b1011000: c <= 9'b111100001;
				8'b101110: c <= 9'b1100100;
				8'b1000001: c <= 9'b10101011;
				default: c <= 9'b0;
			endcase
			9'b10001001 : case(di)
				8'b1000011: c <= 9'b110010100;
				8'b101000: c <= 9'b101111010;
				8'b111010: c <= 9'b110111011;
				8'b110110: c <= 9'b101110001;
				8'b1100100: c <= 9'b110011111;
				8'b1000000: c <= 9'b111010010;
				8'b1110110: c <= 9'b1101111;
				8'b100101: c <= 9'b100011100;
				8'b101111: c <= 9'b111010;
				8'b100110: c <= 9'b100010000;
				8'b1100011: c <= 9'b1100100;
				8'b1001000: c <= 9'b10000;
				8'b111000: c <= 9'b1110111;
				8'b110001: c <= 9'b1100100;
				8'b1010111: c <= 9'b110100;
				8'b1001110: c <= 9'b1111000;
				8'b1101010: c <= 9'b111111110;
				8'b1001001: c <= 9'b1100000;
				8'b1100000: c <= 9'b100100010;
				8'b110111: c <= 9'b100100110;
				8'b1011101: c <= 9'b10001100;
				8'b1011011: c <= 9'b101110101;
				8'b111001: c <= 9'b10111100;
				8'b1001010: c <= 9'b10010001;
				8'b110011: c <= 9'b101100;
				8'b1101100: c <= 9'b1010101;
				8'b1110111: c <= 9'b1101010;
				8'b101011: c <= 9'b111011101;
				8'b1101011: c <= 9'b100010001;
				8'b111100: c <= 9'b110010001;
				8'b1000111: c <= 9'b10000011;
				8'b1011111: c <= 9'b100011000;
				8'b1110100: c <= 9'b10010101;
				8'b101101: c <= 9'b10111011;
				8'b1010011: c <= 9'b110100010;
				8'b1100001: c <= 9'b110001;
				8'b110101: c <= 9'b111100111;
				8'b1000100: c <= 9'b111011101;
				8'b1010001: c <= 9'b1001000;
				8'b1010100: c <= 9'b11011001;
				8'b1100110: c <= 9'b101;
				8'b101010: c <= 9'b1101000;
				8'b1011110: c <= 9'b10110;
				8'b1100111: c <= 9'b101000010;
				8'b1011010: c <= 9'b110101001;
				8'b1000010: c <= 9'b111000110;
				8'b111101: c <= 9'b11001110;
				8'b110000: c <= 9'b10100101;
				8'b111110: c <= 9'b10011101;
				8'b1100010: c <= 9'b100110;
				8'b1110000: c <= 9'b101100000;
				8'b1101001: c <= 9'b1000100;
				8'b1110011: c <= 9'b110;
				8'b1001100: c <= 9'b110011000;
				8'b100001: c <= 9'b100101101;
				8'b1000110: c <= 9'b11100001;
				8'b1110010: c <= 9'b100010000;
				8'b1010000: c <= 9'b1010000;
				8'b1111010: c <= 9'b100011001;
				8'b1010101: c <= 9'b101100010;
				8'b111011: c <= 9'b1011;
				8'b1001101: c <= 9'b100100011;
				8'b111111: c <= 9'b1100111;
				8'b1101110: c <= 9'b11110111;
				8'b1111011: c <= 9'b111001001;
				8'b1001011: c <= 9'b1011001;
				8'b1101111: c <= 9'b1010001;
				8'b1101000: c <= 9'b100011000;
				8'b101100: c <= 9'b1111111;
				8'b100100: c <= 9'b1001110;
				8'b1111000: c <= 9'b101110011;
				8'b1000101: c <= 9'b111000011;
				8'b1011001: c <= 9'b1010101;
				8'b110100: c <= 9'b1010000;
				8'b1111001: c <= 9'b1101100;
				8'b1110001: c <= 9'b1111011;
				8'b1001111: c <= 9'b110000111;
				8'b1100101: c <= 9'b110011000;
				8'b1111110: c <= 9'b10100010;
				8'b1111100: c <= 9'b11000001;
				8'b1010110: c <= 9'b111111001;
				8'b110010: c <= 9'b111011111;
				8'b1101101: c <= 9'b11011100;
				8'b100011: c <= 9'b100101110;
				8'b1110101: c <= 9'b10010011;
				8'b1111101: c <= 9'b10100011;
				8'b101001: c <= 9'b100000000;
				8'b1010010: c <= 9'b101001001;
				8'b1011000: c <= 9'b11100010;
				8'b101110: c <= 9'b111101001;
				8'b1000001: c <= 9'b11101000;
				default: c <= 9'b0;
			endcase
			9'b10011 : case(di)
				8'b1000011: c <= 9'b111110001;
				8'b101000: c <= 9'b100001100;
				8'b111010: c <= 9'b11011110;
				8'b110110: c <= 9'b111010001;
				8'b1100100: c <= 9'b11101001;
				8'b1000000: c <= 9'b111001111;
				8'b1110110: c <= 9'b101010101;
				8'b100101: c <= 9'b110110010;
				8'b101111: c <= 9'b1010111;
				8'b100110: c <= 9'b10100100;
				8'b1100011: c <= 9'b100010000;
				8'b1001000: c <= 9'b101111111;
				8'b111000: c <= 9'b110101;
				8'b110001: c <= 9'b111100;
				8'b1010111: c <= 9'b1110111;
				8'b1001110: c <= 9'b101001111;
				8'b1101010: c <= 9'b1101100;
				8'b1001001: c <= 9'b111111;
				8'b1100000: c <= 9'b101101100;
				8'b110111: c <= 9'b101;
				8'b1011101: c <= 9'b100001111;
				8'b1011011: c <= 9'b1010010;
				8'b111001: c <= 9'b10111000;
				8'b1001010: c <= 9'b11101001;
				8'b110011: c <= 9'b111101001;
				8'b1101100: c <= 9'b100111011;
				8'b1110111: c <= 9'b11100101;
				8'b101011: c <= 9'b101100110;
				8'b1101011: c <= 9'b111100011;
				8'b111100: c <= 9'b110101110;
				8'b1000111: c <= 9'b1101;
				8'b1011111: c <= 9'b10001111;
				8'b1110100: c <= 9'b100;
				8'b101101: c <= 9'b11000100;
				8'b1010011: c <= 9'b100101000;
				8'b1100001: c <= 9'b100010010;
				8'b110101: c <= 9'b111010;
				8'b1000100: c <= 9'b1011000;
				8'b1010001: c <= 9'b11010;
				8'b1010100: c <= 9'b1001011;
				8'b1100110: c <= 9'b11001110;
				8'b101010: c <= 9'b101010111;
				8'b1011110: c <= 9'b111110110;
				8'b1100111: c <= 9'b1100010;
				8'b1011010: c <= 9'b110110000;
				8'b1000010: c <= 9'b101101001;
				8'b111101: c <= 9'b100010100;
				8'b110000: c <= 9'b101101001;
				8'b111110: c <= 9'b101111000;
				8'b1100010: c <= 9'b10101110;
				8'b1110000: c <= 9'b11101001;
				8'b1101001: c <= 9'b11111001;
				8'b1110011: c <= 9'b111101110;
				8'b1001100: c <= 9'b1001010;
				8'b100001: c <= 9'b1110001;
				8'b1000110: c <= 9'b10000011;
				8'b1110010: c <= 9'b110111001;
				8'b1010000: c <= 9'b11111011;
				8'b1111010: c <= 9'b111001111;
				8'b1010101: c <= 9'b111010001;
				8'b111011: c <= 9'b101011011;
				8'b1001101: c <= 9'b101110;
				8'b111111: c <= 9'b10110011;
				8'b1101110: c <= 9'b111110011;
				8'b1111011: c <= 9'b1000111;
				8'b1001011: c <= 9'b100010111;
				8'b1101111: c <= 9'b111111110;
				8'b1101000: c <= 9'b1101010;
				8'b101100: c <= 9'b111010100;
				8'b100100: c <= 9'b1000;
				8'b1111000: c <= 9'b100111110;
				8'b1000101: c <= 9'b110010100;
				8'b1011001: c <= 9'b101100111;
				8'b110100: c <= 9'b1001011;
				8'b1111001: c <= 9'b100100000;
				8'b1110001: c <= 9'b11001;
				8'b1001111: c <= 9'b111111000;
				8'b1100101: c <= 9'b100000001;
				8'b1111110: c <= 9'b101010011;
				8'b1111100: c <= 9'b101;
				8'b1010110: c <= 9'b100011100;
				8'b110010: c <= 9'b111101000;
				8'b1101101: c <= 9'b1010010;
				8'b100011: c <= 9'b100101101;
				8'b1110101: c <= 9'b101100;
				8'b1111101: c <= 9'b111000010;
				8'b101001: c <= 9'b100000101;
				8'b1010010: c <= 9'b10111011;
				8'b1011000: c <= 9'b101111111;
				8'b101110: c <= 9'b111010100;
				8'b1000001: c <= 9'b11101111;
				default: c <= 9'b0;
			endcase
			9'b100101101 : case(di)
				8'b1000011: c <= 9'b1000010;
				8'b101000: c <= 9'b101001110;
				8'b111010: c <= 9'b100000011;
				8'b110110: c <= 9'b11010;
				8'b1100100: c <= 9'b10100000;
				8'b1000000: c <= 9'b100100010;
				8'b1110110: c <= 9'b100110101;
				8'b100101: c <= 9'b111010111;
				8'b101111: c <= 9'b11001110;
				8'b100110: c <= 9'b110011000;
				8'b1100011: c <= 9'b110110111;
				8'b1001000: c <= 9'b101100100;
				8'b111000: c <= 9'b1;
				8'b110001: c <= 9'b10111101;
				8'b1010111: c <= 9'b100001010;
				8'b1001110: c <= 9'b101010010;
				8'b1101010: c <= 9'b110101001;
				8'b1001001: c <= 9'b1011001;
				8'b1100000: c <= 9'b10000101;
				8'b110111: c <= 9'b10101001;
				8'b1011101: c <= 9'b11000010;
				8'b1011011: c <= 9'b10001110;
				8'b111001: c <= 9'b100000100;
				8'b1001010: c <= 9'b111000111;
				8'b110011: c <= 9'b11000110;
				8'b1101100: c <= 9'b1000;
				8'b1110111: c <= 9'b111001100;
				8'b101011: c <= 9'b110100010;
				8'b1101011: c <= 9'b10100;
				8'b111100: c <= 9'b11110;
				8'b1000111: c <= 9'b10110110;
				8'b1011111: c <= 9'b101010001;
				8'b1110100: c <= 9'b101011011;
				8'b101101: c <= 9'b110000;
				8'b1010011: c <= 9'b1001110;
				8'b1100001: c <= 9'b111001101;
				8'b110101: c <= 9'b11000111;
				8'b1000100: c <= 9'b110010010;
				8'b1010001: c <= 9'b10100111;
				8'b1010100: c <= 9'b1000111;
				8'b1100110: c <= 9'b110100000;
				8'b101010: c <= 9'b101000101;
				8'b1011110: c <= 9'b101101001;
				8'b1100111: c <= 9'b101110111;
				8'b1011010: c <= 9'b101010101;
				8'b1000010: c <= 9'b10111011;
				8'b111101: c <= 9'b101110100;
				8'b110000: c <= 9'b10101011;
				8'b111110: c <= 9'b111100001;
				8'b1100010: c <= 9'b10010110;
				8'b1110000: c <= 9'b101010110;
				8'b1101001: c <= 9'b100011011;
				8'b1110011: c <= 9'b10000111;
				8'b1001100: c <= 9'b10100;
				8'b100001: c <= 9'b1111001;
				8'b1000110: c <= 9'b100000111;
				8'b1110010: c <= 9'b10110111;
				8'b1010000: c <= 9'b11110001;
				8'b1111010: c <= 9'b11100101;
				8'b1010101: c <= 9'b111011001;
				8'b111011: c <= 9'b101100100;
				8'b1001101: c <= 9'b11010011;
				8'b111111: c <= 9'b10010101;
				8'b1101110: c <= 9'b1111000;
				8'b1111011: c <= 9'b111001010;
				8'b1001011: c <= 9'b1110011;
				8'b1101111: c <= 9'b1110011;
				8'b1101000: c <= 9'b111110001;
				8'b101100: c <= 9'b111100010;
				8'b100100: c <= 9'b10000010;
				8'b1111000: c <= 9'b10011001;
				8'b1000101: c <= 9'b110000001;
				8'b1011001: c <= 9'b10110001;
				8'b110100: c <= 9'b110100111;
				8'b1111001: c <= 9'b11;
				8'b1110001: c <= 9'b100010111;
				8'b1001111: c <= 9'b101101;
				8'b1100101: c <= 9'b100000001;
				8'b1111110: c <= 9'b100011100;
				8'b1111100: c <= 9'b100100110;
				8'b1010110: c <= 9'b100011011;
				8'b110010: c <= 9'b111011010;
				8'b1101101: c <= 9'b110011001;
				8'b100011: c <= 9'b11111001;
				8'b1110101: c <= 9'b10000111;
				8'b1111101: c <= 9'b100000000;
				8'b101001: c <= 9'b100000100;
				8'b1010010: c <= 9'b101101101;
				8'b1011000: c <= 9'b11111101;
				8'b101110: c <= 9'b10010110;
				8'b1000001: c <= 9'b1101110;
				default: c <= 9'b0;
			endcase
			9'b101001111 : case(di)
				8'b1000011: c <= 9'b101000;
				8'b101000: c <= 9'b10100101;
				8'b111010: c <= 9'b1001110;
				8'b110110: c <= 9'b110100001;
				8'b1100100: c <= 9'b110011000;
				8'b1000000: c <= 9'b110011001;
				8'b1110110: c <= 9'b101110001;
				8'b100101: c <= 9'b11001111;
				8'b101111: c <= 9'b101101000;
				8'b100110: c <= 9'b110011001;
				8'b1100011: c <= 9'b111011;
				8'b1001000: c <= 9'b11011101;
				8'b111000: c <= 9'b10110001;
				8'b110001: c <= 9'b1100101;
				8'b1010111: c <= 9'b111111110;
				8'b1001110: c <= 9'b101100001;
				8'b1101010: c <= 9'b101011110;
				8'b1001001: c <= 9'b10111001;
				8'b1100000: c <= 9'b111010111;
				8'b110111: c <= 9'b110011100;
				8'b1011101: c <= 9'b100010000;
				8'b1011011: c <= 9'b100111111;
				8'b111001: c <= 9'b111011111;
				8'b1001010: c <= 9'b111000011;
				8'b110011: c <= 9'b101000101;
				8'b1101100: c <= 9'b1101101;
				8'b1110111: c <= 9'b100011000;
				8'b101011: c <= 9'b101110010;
				8'b1101011: c <= 9'b11100011;
				8'b111100: c <= 9'b11010000;
				8'b1000111: c <= 9'b1001111;
				8'b1011111: c <= 9'b110011;
				8'b1110100: c <= 9'b110101101;
				8'b101101: c <= 9'b100110010;
				8'b1010011: c <= 9'b10100110;
				8'b1100001: c <= 9'b101100100;
				8'b110101: c <= 9'b100001011;
				8'b1000100: c <= 9'b101110010;
				8'b1010001: c <= 9'b11011101;
				8'b1010100: c <= 9'b11010011;
				8'b1100110: c <= 9'b1011111;
				8'b101010: c <= 9'b1110010;
				8'b1011110: c <= 9'b11101000;
				8'b1100111: c <= 9'b1110;
				8'b1011010: c <= 9'b10101001;
				8'b1000010: c <= 9'b100001010;
				8'b111101: c <= 9'b11101000;
				8'b110000: c <= 9'b111110110;
				8'b111110: c <= 9'b11110001;
				8'b1100010: c <= 9'b101101001;
				8'b1110000: c <= 9'b110011001;
				8'b1101001: c <= 9'b111010110;
				8'b1110011: c <= 9'b10001000;
				8'b1001100: c <= 9'b111010111;
				8'b100001: c <= 9'b1000010;
				8'b1000110: c <= 9'b1010001;
				8'b1110010: c <= 9'b100000010;
				8'b1010000: c <= 9'b100001100;
				8'b1111010: c <= 9'b101011110;
				8'b1010101: c <= 9'b11111101;
				8'b111011: c <= 9'b11101001;
				8'b1001101: c <= 9'b111110110;
				8'b111111: c <= 9'b110111110;
				8'b1101110: c <= 9'b111000000;
				8'b1111011: c <= 9'b1101001;
				8'b1001011: c <= 9'b11110000;
				8'b1101111: c <= 9'b101011011;
				8'b1101000: c <= 9'b10101100;
				8'b101100: c <= 9'b101000100;
				8'b100100: c <= 9'b10100101;
				8'b1111000: c <= 9'b1111011;
				8'b1000101: c <= 9'b11000;
				8'b1011001: c <= 9'b11110100;
				8'b110100: c <= 9'b1100000;
				8'b1111001: c <= 9'b100100;
				8'b1110001: c <= 9'b11110011;
				8'b1001111: c <= 9'b100110;
				8'b1100101: c <= 9'b101011011;
				8'b1111110: c <= 9'b101110011;
				8'b1111100: c <= 9'b110010101;
				8'b1010110: c <= 9'b110001100;
				8'b110010: c <= 9'b1011001;
				8'b1101101: c <= 9'b110110;
				8'b100011: c <= 9'b1000111;
				8'b1110101: c <= 9'b110100;
				8'b1111101: c <= 9'b111010010;
				8'b101001: c <= 9'b110101101;
				8'b1010010: c <= 9'b111110000;
				8'b1011000: c <= 9'b10100101;
				8'b101110: c <= 9'b101010100;
				8'b1000001: c <= 9'b11011;
				default: c <= 9'b0;
			endcase
			9'b101111111 : case(di)
				8'b1000011: c <= 9'b100011011;
				8'b101000: c <= 9'b10111111;
				8'b111010: c <= 9'b111000111;
				8'b110110: c <= 9'b1111110;
				8'b1100100: c <= 9'b1101110;
				8'b1000000: c <= 9'b110100111;
				8'b1110110: c <= 9'b11000010;
				8'b100101: c <= 9'b10001001;
				8'b101111: c <= 9'b10100011;
				8'b100110: c <= 9'b101010000;
				8'b1100011: c <= 9'b100000110;
				8'b1001000: c <= 9'b101101110;
				8'b111000: c <= 9'b11111001;
				8'b110001: c <= 9'b100010011;
				8'b1010111: c <= 9'b11010000;
				8'b1001110: c <= 9'b101110111;
				8'b1101010: c <= 9'b111001000;
				8'b1001001: c <= 9'b111111000;
				8'b1100000: c <= 9'b10111001;
				8'b110111: c <= 9'b101010101;
				8'b1011101: c <= 9'b11111101;
				8'b1011011: c <= 9'b1101101;
				8'b111001: c <= 9'b111011111;
				8'b1001010: c <= 9'b10;
				8'b110011: c <= 9'b100000111;
				8'b1101100: c <= 9'b111100;
				8'b1110111: c <= 9'b1010001;
				8'b101011: c <= 9'b1110011;
				8'b1101011: c <= 9'b100000011;
				8'b111100: c <= 9'b110010110;
				8'b1000111: c <= 9'b11010111;
				8'b1011111: c <= 9'b101100101;
				8'b1110100: c <= 9'b10000011;
				8'b101101: c <= 9'b110011011;
				8'b1010011: c <= 9'b101111110;
				8'b1100001: c <= 9'b101010000;
				8'b110101: c <= 9'b111011011;
				8'b1000100: c <= 9'b10001110;
				8'b1010001: c <= 9'b11001010;
				8'b1010100: c <= 9'b11001110;
				8'b1100110: c <= 9'b10100010;
				8'b101010: c <= 9'b110111011;
				8'b1011110: c <= 9'b110110101;
				8'b1100111: c <= 9'b1010001;
				8'b1011010: c <= 9'b101010100;
				8'b1000010: c <= 9'b10001000;
				8'b111101: c <= 9'b111;
				8'b110000: c <= 9'b110001;
				8'b111110: c <= 9'b1010011;
				8'b1100010: c <= 9'b100011011;
				8'b1110000: c <= 9'b110011111;
				8'b1101001: c <= 9'b1110001;
				8'b1110011: c <= 9'b1001011;
				8'b1001100: c <= 9'b11011011;
				8'b100001: c <= 9'b101110010;
				8'b1000110: c <= 9'b100110111;
				8'b1110010: c <= 9'b111110011;
				8'b1010000: c <= 9'b11000111;
				8'b1111010: c <= 9'b110001100;
				8'b1010101: c <= 9'b11011;
				8'b111011: c <= 9'b101001100;
				8'b1001101: c <= 9'b10001000;
				8'b111111: c <= 9'b110001001;
				8'b1101110: c <= 9'b110110010;
				8'b1111011: c <= 9'b100010110;
				8'b1001011: c <= 9'b10110100;
				8'b1101111: c <= 9'b10010111;
				8'b1101000: c <= 9'b10100111;
				8'b101100: c <= 9'b110011011;
				8'b100100: c <= 9'b111111000;
				8'b1111000: c <= 9'b10110100;
				8'b1000101: c <= 9'b110101011;
				8'b1011001: c <= 9'b111010010;
				8'b110100: c <= 9'b101001111;
				8'b1111001: c <= 9'b1001000;
				8'b1110001: c <= 9'b10101111;
				8'b1001111: c <= 9'b1101001;
				8'b1100101: c <= 9'b101011010;
				8'b1111110: c <= 9'b100100101;
				8'b1111100: c <= 9'b10100101;
				8'b1010110: c <= 9'b101000101;
				8'b110010: c <= 9'b11100100;
				8'b1101101: c <= 9'b11110010;
				8'b100011: c <= 9'b1100010;
				8'b1110101: c <= 9'b100000101;
				8'b1111101: c <= 9'b11010;
				8'b101001: c <= 9'b10000111;
				8'b1010010: c <= 9'b110111010;
				8'b1011000: c <= 9'b1001101;
				8'b101110: c <= 9'b111001111;
				8'b1000001: c <= 9'b111011011;
				default: c <= 9'b0;
			endcase
			9'b1110100 : case(di)
				8'b1000011: c <= 9'b1011111;
				8'b101000: c <= 9'b110001010;
				8'b111010: c <= 9'b11111;
				8'b110110: c <= 9'b101010111;
				8'b1100100: c <= 9'b1111011;
				8'b1000000: c <= 9'b110011010;
				8'b1110110: c <= 9'b111010100;
				8'b100101: c <= 9'b111011100;
				8'b101111: c <= 9'b10101;
				8'b100110: c <= 9'b100101010;
				8'b1100011: c <= 9'b110011001;
				8'b1001000: c <= 9'b100011000;
				8'b111000: c <= 9'b100100001;
				8'b110001: c <= 9'b100101110;
				8'b1010111: c <= 9'b11011100;
				8'b1001110: c <= 9'b110100101;
				8'b1101010: c <= 9'b1111010;
				8'b1001001: c <= 9'b110110100;
				8'b1100000: c <= 9'b100100000;
				8'b110111: c <= 9'b110011001;
				8'b1011101: c <= 9'b101101010;
				8'b1011011: c <= 9'b11101001;
				8'b111001: c <= 9'b11110000;
				8'b1001010: c <= 9'b101010110;
				8'b110011: c <= 9'b110110000;
				8'b1101100: c <= 9'b10011101;
				8'b1110111: c <= 9'b101011011;
				8'b101011: c <= 9'b110111110;
				8'b1101011: c <= 9'b10001100;
				8'b111100: c <= 9'b10100110;
				8'b1000111: c <= 9'b100001101;
				8'b1011111: c <= 9'b11011001;
				8'b1110100: c <= 9'b1010000;
				8'b101101: c <= 9'b110001000;
				8'b1010011: c <= 9'b11001011;
				8'b1100001: c <= 9'b101101001;
				8'b110101: c <= 9'b1000100;
				8'b1000100: c <= 9'b100110111;
				8'b1010001: c <= 9'b101100000;
				8'b1010100: c <= 9'b111111111;
				8'b1100110: c <= 9'b110100001;
				8'b101010: c <= 9'b111101010;
				8'b1011110: c <= 9'b111101110;
				8'b1100111: c <= 9'b100111111;
				8'b1011010: c <= 9'b101110101;
				8'b1000010: c <= 9'b10000111;
				8'b111101: c <= 9'b10010101;
				8'b110000: c <= 9'b101011101;
				8'b111110: c <= 9'b101111010;
				8'b1100010: c <= 9'b110010;
				8'b1110000: c <= 9'b111000110;
				8'b1101001: c <= 9'b1110010;
				8'b1110011: c <= 9'b110100101;
				8'b1001100: c <= 9'b110101011;
				8'b100001: c <= 9'b101101;
				8'b1000110: c <= 9'b111010000;
				8'b1110010: c <= 9'b100011100;
				8'b1010000: c <= 9'b10101111;
				8'b1111010: c <= 9'b11111;
				8'b1010101: c <= 9'b111101110;
				8'b111011: c <= 9'b101011010;
				8'b1001101: c <= 9'b100111101;
				8'b111111: c <= 9'b10010100;
				8'b1101110: c <= 9'b111001;
				8'b1111011: c <= 9'b11000111;
				8'b1001011: c <= 9'b11000010;
				8'b1101111: c <= 9'b100001;
				8'b1101000: c <= 9'b10101101;
				8'b101100: c <= 9'b11;
				8'b100100: c <= 9'b101001000;
				8'b1111000: c <= 9'b1011000;
				8'b1000101: c <= 9'b101110;
				8'b1011001: c <= 9'b101000011;
				8'b110100: c <= 9'b101010001;
				8'b1111001: c <= 9'b110110010;
				8'b1110001: c <= 9'b100000011;
				8'b1001111: c <= 9'b101111110;
				8'b1100101: c <= 9'b111;
				8'b1111110: c <= 9'b10101110;
				8'b1111100: c <= 9'b111111101;
				8'b1010110: c <= 9'b11101000;
				8'b110010: c <= 9'b1100010;
				8'b1101101: c <= 9'b100110010;
				8'b100011: c <= 9'b110010;
				8'b1110101: c <= 9'b100011;
				8'b1111101: c <= 9'b100100001;
				8'b101001: c <= 9'b111100111;
				8'b1010010: c <= 9'b111101111;
				8'b1011000: c <= 9'b11110000;
				8'b101110: c <= 9'b10011;
				8'b1000001: c <= 9'b111010100;
				default: c <= 9'b0;
			endcase
			9'b110000 : case(di)
				8'b1000011: c <= 9'b11111101;
				8'b101000: c <= 9'b101100;
				8'b111010: c <= 9'b101011101;
				8'b110110: c <= 9'b101001011;
				8'b1100100: c <= 9'b111000010;
				8'b1000000: c <= 9'b101000100;
				8'b1110110: c <= 9'b101001010;
				8'b100101: c <= 9'b100011001;
				8'b101111: c <= 9'b101010100;
				8'b100110: c <= 9'b100001;
				8'b1100011: c <= 9'b11100101;
				8'b1001000: c <= 9'b110000001;
				8'b111000: c <= 9'b10100011;
				8'b110001: c <= 9'b11011000;
				8'b1010111: c <= 9'b111000110;
				8'b1001110: c <= 9'b111011110;
				8'b1101010: c <= 9'b100001111;
				8'b1001001: c <= 9'b10101011;
				8'b1100000: c <= 9'b10011100;
				8'b110111: c <= 9'b10101101;
				8'b1011101: c <= 9'b10100111;
				8'b1011011: c <= 9'b110101111;
				8'b111001: c <= 9'b100010010;
				8'b1001010: c <= 9'b110011111;
				8'b110011: c <= 9'b1;
				8'b1101100: c <= 9'b100010000;
				8'b1110111: c <= 9'b11011101;
				8'b101011: c <= 9'b1000111;
				8'b1101011: c <= 9'b1110001;
				8'b111100: c <= 9'b101011;
				8'b1000111: c <= 9'b10100000;
				8'b1011111: c <= 9'b1;
				8'b1110100: c <= 9'b10101011;
				8'b101101: c <= 9'b1011110;
				8'b1010011: c <= 9'b1111010;
				8'b1100001: c <= 9'b110000000;
				8'b110101: c <= 9'b10110010;
				8'b1000100: c <= 9'b10110111;
				8'b1010001: c <= 9'b100001101;
				8'b1010100: c <= 9'b101011001;
				8'b1100110: c <= 9'b111011;
				8'b101010: c <= 9'b100011011;
				8'b1011110: c <= 9'b111001101;
				8'b1100111: c <= 9'b100100010;
				8'b1011010: c <= 9'b111110001;
				8'b1000010: c <= 9'b10111010;
				8'b111101: c <= 9'b100010000;
				8'b110000: c <= 9'b10100111;
				8'b111110: c <= 9'b111111101;
				8'b1100010: c <= 9'b100001111;
				8'b1110000: c <= 9'b100001111;
				8'b1101001: c <= 9'b110101011;
				8'b1110011: c <= 9'b11100001;
				8'b1001100: c <= 9'b100000000;
				8'b100001: c <= 9'b100011000;
				8'b1000110: c <= 9'b100001101;
				8'b1110010: c <= 9'b10100;
				8'b1010000: c <= 9'b10010100;
				8'b1111010: c <= 9'b1011100;
				8'b1010101: c <= 9'b100101011;
				8'b111011: c <= 9'b101011;
				8'b1001101: c <= 9'b1111110;
				8'b111111: c <= 9'b10101010;
				8'b1101110: c <= 9'b100100000;
				8'b1111011: c <= 9'b111000000;
				8'b1001011: c <= 9'b101011010;
				8'b1101111: c <= 9'b10101101;
				8'b1101000: c <= 9'b101010100;
				8'b101100: c <= 9'b101000010;
				8'b100100: c <= 9'b10001010;
				8'b1111000: c <= 9'b10111100;
				8'b1000101: c <= 9'b110000001;
				8'b1011001: c <= 9'b100110100;
				8'b110100: c <= 9'b110111000;
				8'b1111001: c <= 9'b11001100;
				8'b1110001: c <= 9'b110011010;
				8'b1001111: c <= 9'b11100111;
				8'b1100101: c <= 9'b101101100;
				8'b1111110: c <= 9'b110000110;
				8'b1111100: c <= 9'b110010001;
				8'b1010110: c <= 9'b100001110;
				8'b110010: c <= 9'b11110110;
				8'b1101101: c <= 9'b110001000;
				8'b100011: c <= 9'b1111010;
				8'b1110101: c <= 9'b111011111;
				8'b1111101: c <= 9'b11110111;
				8'b101001: c <= 9'b1010000;
				8'b1010010: c <= 9'b1001111;
				8'b1011000: c <= 9'b101101;
				8'b101110: c <= 9'b100011010;
				8'b1000001: c <= 9'b11001111;
				default: c <= 9'b0;
			endcase
			9'b1001010 : case(di)
				8'b1000011: c <= 9'b110111001;
				8'b101000: c <= 9'b10000000;
				8'b111010: c <= 9'b111111011;
				8'b110110: c <= 9'b10001011;
				8'b1100100: c <= 9'b1101;
				8'b1000000: c <= 9'b100001011;
				8'b1110110: c <= 9'b101000110;
				8'b100101: c <= 9'b110110101;
				8'b101111: c <= 9'b110110011;
				8'b100110: c <= 9'b11110011;
				8'b1100011: c <= 9'b101010110;
				8'b1001000: c <= 9'b100100111;
				8'b111000: c <= 9'b111111;
				8'b110001: c <= 9'b10011000;
				8'b1010111: c <= 9'b10101;
				8'b1001110: c <= 9'b110100100;
				8'b1101010: c <= 9'b101110010;
				8'b1001001: c <= 9'b100001001;
				8'b1100000: c <= 9'b11101111;
				8'b110111: c <= 9'b111011110;
				8'b1011101: c <= 9'b1010111;
				8'b1011011: c <= 9'b100110111;
				8'b111001: c <= 9'b1000100;
				8'b1001010: c <= 9'b11011100;
				8'b110011: c <= 9'b1101010;
				8'b1101100: c <= 9'b1110011;
				8'b1110111: c <= 9'b100001111;
				8'b101011: c <= 9'b100001111;
				8'b1101011: c <= 9'b11011001;
				8'b111100: c <= 9'b111000010;
				8'b1000111: c <= 9'b10100111;
				8'b1011111: c <= 9'b10110011;
				8'b1110100: c <= 9'b111000110;
				8'b101101: c <= 9'b101100001;
				8'b1010011: c <= 9'b10101100;
				8'b1100001: c <= 9'b110000001;
				8'b110101: c <= 9'b100000101;
				8'b1000100: c <= 9'b100110100;
				8'b1010001: c <= 9'b111001001;
				8'b1010100: c <= 9'b100001;
				8'b1100110: c <= 9'b110101111;
				8'b101010: c <= 9'b110111011;
				8'b1011110: c <= 9'b110101110;
				8'b1100111: c <= 9'b1100100;
				8'b1011010: c <= 9'b11101000;
				8'b1000010: c <= 9'b110001110;
				8'b111101: c <= 9'b11011010;
				8'b110000: c <= 9'b100111011;
				8'b111110: c <= 9'b11010010;
				8'b1100010: c <= 9'b101010010;
				8'b1110000: c <= 9'b1001010;
				8'b1101001: c <= 9'b101110001;
				8'b1110011: c <= 9'b111110011;
				8'b1001100: c <= 9'b1111101;
				8'b100001: c <= 9'b101011110;
				8'b1000110: c <= 9'b11000;
				8'b1110010: c <= 9'b100100010;
				8'b1010000: c <= 9'b101101000;
				8'b1111010: c <= 9'b100011111;
				8'b1010101: c <= 9'b100010001;
				8'b111011: c <= 9'b1100110;
				8'b1001101: c <= 9'b1110111;
				8'b111111: c <= 9'b110011000;
				8'b1101110: c <= 9'b111000;
				8'b1111011: c <= 9'b110000010;
				8'b1001011: c <= 9'b111101000;
				8'b1101111: c <= 9'b100010101;
				8'b1101000: c <= 9'b10110111;
				8'b101100: c <= 9'b11100001;
				8'b100100: c <= 9'b100101110;
				8'b1111000: c <= 9'b101011;
				8'b1000101: c <= 9'b100010;
				8'b1011001: c <= 9'b101010001;
				8'b110100: c <= 9'b111111010;
				8'b1111001: c <= 9'b11111010;
				8'b1110001: c <= 9'b111100101;
				8'b1001111: c <= 9'b100101111;
				8'b1100101: c <= 9'b11010000;
				8'b1111110: c <= 9'b11100111;
				8'b1111100: c <= 9'b101101000;
				8'b1010110: c <= 9'b10011100;
				8'b110010: c <= 9'b100011001;
				8'b1101101: c <= 9'b10000;
				8'b100011: c <= 9'b111111;
				8'b1110101: c <= 9'b10100100;
				8'b1111101: c <= 9'b110001010;
				8'b101001: c <= 9'b110001010;
				8'b1010010: c <= 9'b110011;
				8'b1011000: c <= 9'b1100;
				8'b101110: c <= 9'b110111111;
				8'b1000001: c <= 9'b1001101;
				default: c <= 9'b0;
			endcase
			9'b110010011 : case(di)
				8'b1000011: c <= 9'b10100000;
				8'b101000: c <= 9'b101110111;
				8'b111010: c <= 9'b101110011;
				8'b110110: c <= 9'b101010101;
				8'b1100100: c <= 9'b101111111;
				8'b1000000: c <= 9'b100100011;
				8'b1110110: c <= 9'b111010100;
				8'b100101: c <= 9'b11110100;
				8'b101111: c <= 9'b1000111;
				8'b100110: c <= 9'b11100000;
				8'b1100011: c <= 9'b1010101;
				8'b1001000: c <= 9'b100100010;
				8'b111000: c <= 9'b11101100;
				8'b110001: c <= 9'b11001101;
				8'b1010111: c <= 9'b111101001;
				8'b1001110: c <= 9'b101101111;
				8'b1101010: c <= 9'b111111101;
				8'b1001001: c <= 9'b11100001;
				8'b1100000: c <= 9'b100111001;
				8'b110111: c <= 9'b101000001;
				8'b1011101: c <= 9'b1110001;
				8'b1011011: c <= 9'b10101001;
				8'b111001: c <= 9'b10111000;
				8'b1001010: c <= 9'b100110010;
				8'b110011: c <= 9'b10010110;
				8'b1101100: c <= 9'b10001001;
				8'b1110111: c <= 9'b1100101;
				8'b101011: c <= 9'b101100010;
				8'b1101011: c <= 9'b101101100;
				8'b111100: c <= 9'b10;
				8'b1000111: c <= 9'b10111010;
				8'b1011111: c <= 9'b110100000;
				8'b1110100: c <= 9'b1110100;
				8'b101101: c <= 9'b100101000;
				8'b1010011: c <= 9'b10110011;
				8'b1100001: c <= 9'b10100;
				8'b110101: c <= 9'b10110011;
				8'b1000100: c <= 9'b1011000;
				8'b1010001: c <= 9'b110111000;
				8'b1010100: c <= 9'b110010100;
				8'b1100110: c <= 9'b110000;
				8'b101010: c <= 9'b1100110;
				8'b1011110: c <= 9'b100110110;
				8'b1100111: c <= 9'b1011000;
				8'b1011010: c <= 9'b111010100;
				8'b1000010: c <= 9'b11110111;
				8'b111101: c <= 9'b100011000;
				8'b110000: c <= 9'b110001000;
				8'b111110: c <= 9'b1111001;
				8'b1100010: c <= 9'b11100010;
				8'b1110000: c <= 9'b11110100;
				8'b1101001: c <= 9'b11011011;
				8'b1110011: c <= 9'b101001;
				8'b1001100: c <= 9'b1001111;
				8'b100001: c <= 9'b101011001;
				8'b1000110: c <= 9'b11110;
				8'b1110010: c <= 9'b10111111;
				8'b1010000: c <= 9'b10101;
				8'b1111010: c <= 9'b110001011;
				8'b1010101: c <= 9'b110100101;
				8'b111011: c <= 9'b1000;
				8'b1001101: c <= 9'b11110110;
				8'b111111: c <= 9'b10101010;
				8'b1101110: c <= 9'b1101100;
				8'b1111011: c <= 9'b11111110;
				8'b1001011: c <= 9'b1000000;
				8'b1101111: c <= 9'b110001001;
				8'b1101000: c <= 9'b110100000;
				8'b101100: c <= 9'b100011011;
				8'b100100: c <= 9'b1000011;
				8'b1111000: c <= 9'b101110;
				8'b1000101: c <= 9'b111101010;
				8'b1011001: c <= 9'b1011110;
				8'b110100: c <= 9'b1001001;
				8'b1111001: c <= 9'b10001110;
				8'b1110001: c <= 9'b10000000;
				8'b1001111: c <= 9'b101100100;
				8'b1100101: c <= 9'b110110;
				8'b1111110: c <= 9'b101100011;
				8'b1111100: c <= 9'b11011110;
				8'b1010110: c <= 9'b111011001;
				8'b110010: c <= 9'b111100;
				8'b1101101: c <= 9'b100111110;
				8'b100011: c <= 9'b10110111;
				8'b1110101: c <= 9'b1100110;
				8'b1111101: c <= 9'b101111001;
				8'b101001: c <= 9'b10010100;
				8'b1010010: c <= 9'b111101101;
				8'b1011000: c <= 9'b1100010;
				8'b101110: c <= 9'b100001001;
				8'b1000001: c <= 9'b101110001;
				default: c <= 9'b0;
			endcase
			9'b110111011 : case(di)
				8'b1000011: c <= 9'b1111001;
				8'b101000: c <= 9'b110101111;
				8'b111010: c <= 9'b110110011;
				8'b110110: c <= 9'b100010;
				8'b1100100: c <= 9'b10000010;
				8'b1000000: c <= 9'b111100001;
				8'b1110110: c <= 9'b100111011;
				8'b100101: c <= 9'b111110110;
				8'b101111: c <= 9'b110100010;
				8'b100110: c <= 9'b1111;
				8'b1100011: c <= 9'b10010111;
				8'b1001000: c <= 9'b111100000;
				8'b111000: c <= 9'b1111011;
				8'b110001: c <= 9'b110011110;
				8'b1010111: c <= 9'b100101100;
				8'b1001110: c <= 9'b111001011;
				8'b1101010: c <= 9'b111100101;
				8'b1001001: c <= 9'b10111001;
				8'b1100000: c <= 9'b1110101;
				8'b110111: c <= 9'b10001001;
				8'b1011101: c <= 9'b100011010;
				8'b1011011: c <= 9'b110001100;
				8'b111001: c <= 9'b111001011;
				8'b1001010: c <= 9'b100101011;
				8'b110011: c <= 9'b111010001;
				8'b1101100: c <= 9'b10010100;
				8'b1110111: c <= 9'b1111000;
				8'b101011: c <= 9'b110110;
				8'b1101011: c <= 9'b11101011;
				8'b111100: c <= 9'b101010000;
				8'b1000111: c <= 9'b110000001;
				8'b1011111: c <= 9'b10001110;
				8'b1110100: c <= 9'b1111110;
				8'b101101: c <= 9'b100110010;
				8'b1010011: c <= 9'b101011110;
				8'b1100001: c <= 9'b10111000;
				8'b110101: c <= 9'b10111100;
				8'b1000100: c <= 9'b110;
				8'b1010001: c <= 9'b111010111;
				8'b1010100: c <= 9'b111;
				8'b1100110: c <= 9'b111000011;
				8'b101010: c <= 9'b101010010;
				8'b1011110: c <= 9'b111101110;
				8'b1100111: c <= 9'b10111110;
				8'b1011010: c <= 9'b11010011;
				8'b1000010: c <= 9'b100110000;
				8'b111101: c <= 9'b1111100;
				8'b110000: c <= 9'b110010100;
				8'b111110: c <= 9'b100011100;
				8'b1100010: c <= 9'b110110110;
				8'b1110000: c <= 9'b100;
				8'b1101001: c <= 9'b10011010;
				8'b1110011: c <= 9'b111101001;
				8'b1001100: c <= 9'b10000001;
				8'b100001: c <= 9'b10010011;
				8'b1000110: c <= 9'b101001110;
				8'b1110010: c <= 9'b1101111;
				8'b1010000: c <= 9'b11000011;
				8'b1111010: c <= 9'b1100001;
				8'b1010101: c <= 9'b1101101;
				8'b111011: c <= 9'b111000;
				8'b1001101: c <= 9'b101011101;
				8'b111111: c <= 9'b1011011;
				8'b1101110: c <= 9'b1001100;
				8'b1111011: c <= 9'b10011;
				8'b1001011: c <= 9'b110011000;
				8'b1101111: c <= 9'b10001001;
				8'b1101000: c <= 9'b1000001;
				8'b101100: c <= 9'b110110111;
				8'b100100: c <= 9'b11111100;
				8'b1111000: c <= 9'b11110100;
				8'b1000101: c <= 9'b1011111;
				8'b1011001: c <= 9'b10010011;
				8'b110100: c <= 9'b1100011;
				8'b1111001: c <= 9'b111011111;
				8'b1110001: c <= 9'b10000010;
				8'b1001111: c <= 9'b101100110;
				8'b1100101: c <= 9'b101011;
				8'b1111110: c <= 9'b1000100;
				8'b1111100: c <= 9'b101001010;
				8'b1010110: c <= 9'b1110;
				8'b110010: c <= 9'b111010100;
				8'b1101101: c <= 9'b101010111;
				8'b100011: c <= 9'b111000101;
				8'b1110101: c <= 9'b10101;
				8'b1111101: c <= 9'b11110000;
				8'b101001: c <= 9'b10110011;
				8'b1010010: c <= 9'b110111010;
				8'b1011000: c <= 9'b1101110;
				8'b101110: c <= 9'b11111011;
				8'b1000001: c <= 9'b101100;
				default: c <= 9'b0;
			endcase
			9'b100010 : case(di)
				8'b1000011: c <= 9'b10100110;
				8'b101000: c <= 9'b10000011;
				8'b111010: c <= 9'b110001110;
				8'b110110: c <= 9'b10100000;
				8'b1100100: c <= 9'b111001100;
				8'b1000000: c <= 9'b10000001;
				8'b1110110: c <= 9'b11100101;
				8'b100101: c <= 9'b11011000;
				8'b101111: c <= 9'b100000000;
				8'b100110: c <= 9'b110;
				8'b1100011: c <= 9'b101100110;
				8'b1001000: c <= 9'b110011010;
				8'b111000: c <= 9'b110001;
				8'b110001: c <= 9'b111011100;
				8'b1010111: c <= 9'b1100011;
				8'b1001110: c <= 9'b111111101;
				8'b1101010: c <= 9'b101000001;
				8'b1001001: c <= 9'b1010001;
				8'b1100000: c <= 9'b11110011;
				8'b110111: c <= 9'b10000011;
				8'b1011101: c <= 9'b10111110;
				8'b1011011: c <= 9'b10101100;
				8'b111001: c <= 9'b100011100;
				8'b1001010: c <= 9'b11010101;
				8'b110011: c <= 9'b111100110;
				8'b1101100: c <= 9'b101101011;
				8'b1110111: c <= 9'b110000000;
				8'b101011: c <= 9'b111111001;
				8'b1101011: c <= 9'b110001100;
				8'b111100: c <= 9'b111010010;
				8'b1000111: c <= 9'b110001010;
				8'b1011111: c <= 9'b100101101;
				8'b1110100: c <= 9'b110100001;
				8'b101101: c <= 9'b101001001;
				8'b1010011: c <= 9'b11101011;
				8'b1100001: c <= 9'b111011101;
				8'b110101: c <= 9'b11000110;
				8'b1000100: c <= 9'b100111011;
				8'b1010001: c <= 9'b101000011;
				8'b1010100: c <= 9'b10101000;
				8'b1100110: c <= 9'b100001010;
				8'b101010: c <= 9'b110011000;
				8'b1011110: c <= 9'b101111111;
				8'b1100111: c <= 9'b110010001;
				8'b1011010: c <= 9'b100110010;
				8'b1000010: c <= 9'b110001000;
				8'b111101: c <= 9'b10101;
				8'b110000: c <= 9'b110110010;
				8'b111110: c <= 9'b11111000;
				8'b1100010: c <= 9'b101001111;
				8'b1110000: c <= 9'b111111111;
				8'b1101001: c <= 9'b101001011;
				8'b1110011: c <= 9'b1011000;
				8'b1001100: c <= 9'b11000111;
				8'b100001: c <= 9'b10000011;
				8'b1000110: c <= 9'b101000001;
				8'b1110010: c <= 9'b100110010;
				8'b1010000: c <= 9'b100011;
				8'b1111010: c <= 9'b101001000;
				8'b1010101: c <= 9'b101010110;
				8'b111011: c <= 9'b10000011;
				8'b1001101: c <= 9'b110101;
				8'b111111: c <= 9'b101000001;
				8'b1101110: c <= 9'b101101110;
				8'b1111011: c <= 9'b111111101;
				8'b1001011: c <= 9'b11101000;
				8'b1101111: c <= 9'b110011001;
				8'b1101000: c <= 9'b1111100;
				8'b101100: c <= 9'b100010101;
				8'b100100: c <= 9'b11110110;
				8'b1111000: c <= 9'b1011000;
				8'b1000101: c <= 9'b11011000;
				8'b1011001: c <= 9'b101101;
				8'b110100: c <= 9'b11001101;
				8'b1111001: c <= 9'b1010000;
				8'b1110001: c <= 9'b100001110;
				8'b1001111: c <= 9'b110101110;
				8'b1100101: c <= 9'b1010000;
				8'b1111110: c <= 9'b101011010;
				8'b1111100: c <= 9'b111011;
				8'b1010110: c <= 9'b11110101;
				8'b110010: c <= 9'b10110100;
				8'b1101101: c <= 9'b110011101;
				8'b100011: c <= 9'b100010001;
				8'b1110101: c <= 9'b11010;
				8'b1111101: c <= 9'b110000010;
				8'b101001: c <= 9'b11101111;
				8'b1010010: c <= 9'b110110111;
				8'b1011000: c <= 9'b100100000;
				8'b101110: c <= 9'b101101011;
				8'b1000001: c <= 9'b100111110;
				default: c <= 9'b0;
			endcase
			9'b100100101 : case(di)
				8'b1000011: c <= 9'b111011110;
				8'b101000: c <= 9'b1110001;
				8'b111010: c <= 9'b10010100;
				8'b110110: c <= 9'b101101100;
				8'b1100100: c <= 9'b10111110;
				8'b1000000: c <= 9'b11110010;
				8'b1110110: c <= 9'b110010;
				8'b100101: c <= 9'b1000110;
				8'b101111: c <= 9'b1001001;
				8'b100110: c <= 9'b101001000;
				8'b1100011: c <= 9'b101011011;
				8'b1001000: c <= 9'b10111110;
				8'b111000: c <= 9'b100110111;
				8'b110001: c <= 9'b111101010;
				8'b1010111: c <= 9'b101011110;
				8'b1001110: c <= 9'b111101000;
				8'b1101010: c <= 9'b1000111;
				8'b1001001: c <= 9'b10110110;
				8'b1100000: c <= 9'b100010101;
				8'b110111: c <= 9'b10001000;
				8'b1011101: c <= 9'b110010010;
				8'b1011011: c <= 9'b111110101;
				8'b111001: c <= 9'b10011011;
				8'b1001010: c <= 9'b111010111;
				8'b110011: c <= 9'b1110111;
				8'b1101100: c <= 9'b111101000;
				8'b1110111: c <= 9'b10000110;
				8'b101011: c <= 9'b10101100;
				8'b1101011: c <= 9'b100000100;
				8'b111100: c <= 9'b110110010;
				8'b1000111: c <= 9'b110001000;
				8'b1011111: c <= 9'b11110110;
				8'b1110100: c <= 9'b1011001;
				8'b101101: c <= 9'b1100001;
				8'b1010011: c <= 9'b110000011;
				8'b1100001: c <= 9'b111000000;
				8'b110101: c <= 9'b10000011;
				8'b1000100: c <= 9'b111100011;
				8'b1010001: c <= 9'b11001010;
				8'b1010100: c <= 9'b101010110;
				8'b1100110: c <= 9'b110100101;
				8'b101010: c <= 9'b100010;
				8'b1011110: c <= 9'b1110011;
				8'b1100111: c <= 9'b111000010;
				8'b1011010: c <= 9'b100010100;
				8'b1000010: c <= 9'b11110000;
				8'b111101: c <= 9'b111100100;
				8'b110000: c <= 9'b110001011;
				8'b111110: c <= 9'b100010001;
				8'b1100010: c <= 9'b101111010;
				8'b1110000: c <= 9'b101110001;
				8'b1101001: c <= 9'b110001101;
				8'b1110011: c <= 9'b1011;
				8'b1001100: c <= 9'b111010100;
				8'b100001: c <= 9'b110111100;
				8'b1000110: c <= 9'b100101101;
				8'b1110010: c <= 9'b100100000;
				8'b1010000: c <= 9'b1100101;
				8'b1111010: c <= 9'b110100101;
				8'b1010101: c <= 9'b10001001;
				8'b111011: c <= 9'b111011010;
				8'b1001101: c <= 9'b100000101;
				8'b111111: c <= 9'b10101011;
				8'b1101110: c <= 9'b100010000;
				8'b1111011: c <= 9'b111111111;
				8'b1001011: c <= 9'b1101110;
				8'b1101111: c <= 9'b110111;
				8'b1101000: c <= 9'b1000000;
				8'b101100: c <= 9'b11110101;
				8'b100100: c <= 9'b10001001;
				8'b1111000: c <= 9'b10011000;
				8'b1000101: c <= 9'b11110100;
				8'b1011001: c <= 9'b11111100;
				8'b110100: c <= 9'b100111010;
				8'b1111001: c <= 9'b101100;
				8'b1110001: c <= 9'b111111001;
				8'b1001111: c <= 9'b100100011;
				8'b1100101: c <= 9'b110110000;
				8'b1111110: c <= 9'b10100011;
				8'b1111100: c <= 9'b11101101;
				8'b1010110: c <= 9'b10000;
				8'b110010: c <= 9'b111001010;
				8'b1101101: c <= 9'b11111100;
				8'b100011: c <= 9'b111011110;
				8'b1110101: c <= 9'b10010001;
				8'b1111101: c <= 9'b101110101;
				8'b101001: c <= 9'b10110110;
				8'b1010010: c <= 9'b10111000;
				8'b1011000: c <= 9'b100100101;
				8'b101110: c <= 9'b110000;
				8'b1000001: c <= 9'b111111001;
				default: c <= 9'b0;
			endcase
			9'b100001100 : case(di)
				8'b1000011: c <= 9'b11111101;
				8'b101000: c <= 9'b101100011;
				8'b111010: c <= 9'b100100001;
				8'b110110: c <= 9'b110101111;
				8'b1100100: c <= 9'b100111110;
				8'b1000000: c <= 9'b101111000;
				8'b1110110: c <= 9'b111010010;
				8'b100101: c <= 9'b1111011;
				8'b101111: c <= 9'b11000100;
				8'b100110: c <= 9'b100111111;
				8'b1100011: c <= 9'b100111000;
				8'b1001000: c <= 9'b1111111;
				8'b111000: c <= 9'b111111011;
				8'b110001: c <= 9'b10000110;
				8'b1010111: c <= 9'b1111101;
				8'b1001110: c <= 9'b1110;
				8'b1101010: c <= 9'b100110011;
				8'b1001001: c <= 9'b101101101;
				8'b1100000: c <= 9'b110111110;
				8'b110111: c <= 9'b101001011;
				8'b1011101: c <= 9'b110111111;
				8'b1011011: c <= 9'b100011000;
				8'b111001: c <= 9'b10101101;
				8'b1001010: c <= 9'b100001100;
				8'b110011: c <= 9'b1010110;
				8'b1101100: c <= 9'b10111001;
				8'b1110111: c <= 9'b101101100;
				8'b101011: c <= 9'b10101000;
				8'b1101011: c <= 9'b101011001;
				8'b111100: c <= 9'b100101101;
				8'b1000111: c <= 9'b100101111;
				8'b1011111: c <= 9'b11010010;
				8'b1110100: c <= 9'b110110011;
				8'b101101: c <= 9'b10100;
				8'b1010011: c <= 9'b11000111;
				8'b1100001: c <= 9'b101011111;
				8'b110101: c <= 9'b100111;
				8'b1000100: c <= 9'b111100001;
				8'b1010001: c <= 9'b111101111;
				8'b1010100: c <= 9'b101110001;
				8'b1100110: c <= 9'b110101111;
				8'b101010: c <= 9'b1001100;
				8'b1011110: c <= 9'b10001110;
				8'b1100111: c <= 9'b10100111;
				8'b1011010: c <= 9'b11000110;
				8'b1000010: c <= 9'b110011010;
				8'b111101: c <= 9'b111111010;
				8'b110000: c <= 9'b111101101;
				8'b111110: c <= 9'b100000111;
				8'b1100010: c <= 9'b101110010;
				8'b1110000: c <= 9'b11101001;
				8'b1101001: c <= 9'b10011111;
				8'b1110011: c <= 9'b111001100;
				8'b1001100: c <= 9'b100001001;
				8'b100001: c <= 9'b1111111;
				8'b1000110: c <= 9'b111100010;
				8'b1110010: c <= 9'b11110100;
				8'b1010000: c <= 9'b11011010;
				8'b1111010: c <= 9'b111010000;
				8'b1010101: c <= 9'b110000101;
				8'b111011: c <= 9'b100011100;
				8'b1001101: c <= 9'b11110111;
				8'b111111: c <= 9'b101110010;
				8'b1101110: c <= 9'b110110011;
				8'b1111011: c <= 9'b11000011;
				8'b1001011: c <= 9'b100110011;
				8'b1101111: c <= 9'b1101001;
				8'b1101000: c <= 9'b11110011;
				8'b101100: c <= 9'b101001100;
				8'b100100: c <= 9'b100101011;
				8'b1111000: c <= 9'b100110110;
				8'b1000101: c <= 9'b110011;
				8'b1011001: c <= 9'b1100000;
				8'b110100: c <= 9'b10100111;
				8'b1111001: c <= 9'b110011101;
				8'b1110001: c <= 9'b1111001;
				8'b1001111: c <= 9'b10101101;
				8'b1100101: c <= 9'b111110000;
				8'b1111110: c <= 9'b100010000;
				8'b1111100: c <= 9'b100101100;
				8'b1010110: c <= 9'b11100110;
				8'b110010: c <= 9'b111100;
				8'b1101101: c <= 9'b1000;
				8'b100011: c <= 9'b10100101;
				8'b1110101: c <= 9'b111000100;
				8'b1111101: c <= 9'b101101000;
				8'b101001: c <= 9'b100011100;
				8'b1010010: c <= 9'b100000011;
				8'b1011000: c <= 9'b10110;
				8'b101110: c <= 9'b111010;
				8'b1000001: c <= 9'b100001100;
				default: c <= 9'b0;
			endcase
			9'b10011000 : case(di)
				8'b1000011: c <= 9'b10011011;
				8'b101000: c <= 9'b110110010;
				8'b111010: c <= 9'b110001100;
				8'b110110: c <= 9'b110111011;
				8'b1100100: c <= 9'b110100101;
				8'b1000000: c <= 9'b10000011;
				8'b1110110: c <= 9'b110110011;
				8'b100101: c <= 9'b110101011;
				8'b101111: c <= 9'b11000;
				8'b100110: c <= 9'b11101000;
				8'b1100011: c <= 9'b100010100;
				8'b1001000: c <= 9'b100101110;
				8'b111000: c <= 9'b11111110;
				8'b110001: c <= 9'b1101100;
				8'b1010111: c <= 9'b110001000;
				8'b1001110: c <= 9'b1010001;
				8'b1101010: c <= 9'b110001001;
				8'b1001001: c <= 9'b11111010;
				8'b1100000: c <= 9'b10110101;
				8'b110111: c <= 9'b100100111;
				8'b1011101: c <= 9'b101101100;
				8'b1011011: c <= 9'b110011110;
				8'b111001: c <= 9'b11001;
				8'b1001010: c <= 9'b1010001;
				8'b110011: c <= 9'b10100111;
				8'b1101100: c <= 9'b11111101;
				8'b1110111: c <= 9'b10000001;
				8'b101011: c <= 9'b11000111;
				8'b1101011: c <= 9'b100001001;
				8'b111100: c <= 9'b100011011;
				8'b1000111: c <= 9'b101001000;
				8'b1011111: c <= 9'b10001010;
				8'b1110100: c <= 9'b100101111;
				8'b101101: c <= 9'b110010111;
				8'b1010011: c <= 9'b110100001;
				8'b1100001: c <= 9'b111100101;
				8'b110101: c <= 9'b101111110;
				8'b1000100: c <= 9'b11110;
				8'b1010001: c <= 9'b10110110;
				8'b1010100: c <= 9'b111101110;
				8'b1100110: c <= 9'b100010010;
				8'b101010: c <= 9'b101000001;
				8'b1011110: c <= 9'b10010;
				8'b1100111: c <= 9'b100101000;
				8'b1011010: c <= 9'b110001;
				8'b1000010: c <= 9'b10001111;
				8'b111101: c <= 9'b110010011;
				8'b110000: c <= 9'b101010;
				8'b111110: c <= 9'b100111011;
				8'b1100010: c <= 9'b10101100;
				8'b1110000: c <= 9'b100111;
				8'b1101001: c <= 9'b101010011;
				8'b1110011: c <= 9'b101110100;
				8'b1001100: c <= 9'b101000111;
				8'b100001: c <= 9'b101101110;
				8'b1000110: c <= 9'b101100010;
				8'b1110010: c <= 9'b11101000;
				8'b1010000: c <= 9'b11101;
				8'b1111010: c <= 9'b1101001;
				8'b1010101: c <= 9'b111011100;
				8'b111011: c <= 9'b1111001;
				8'b1001101: c <= 9'b101110001;
				8'b111111: c <= 9'b101001000;
				8'b1101110: c <= 9'b110001001;
				8'b1111011: c <= 9'b111111000;
				8'b1001011: c <= 9'b110001101;
				8'b1101111: c <= 9'b1111011;
				8'b1101000: c <= 9'b100011101;
				8'b101100: c <= 9'b10001101;
				8'b100100: c <= 9'b101011111;
				8'b1111000: c <= 9'b11111100;
				8'b1000101: c <= 9'b111100001;
				8'b1011001: c <= 9'b10001011;
				8'b110100: c <= 9'b100010101;
				8'b1111001: c <= 9'b100101010;
				8'b1110001: c <= 9'b1000101;
				8'b1001111: c <= 9'b1110010;
				8'b1100101: c <= 9'b10000101;
				8'b1111110: c <= 9'b10001011;
				8'b1111100: c <= 9'b10011100;
				8'b1010110: c <= 9'b111101101;
				8'b110010: c <= 9'b1111;
				8'b1101101: c <= 9'b101010100;
				8'b100011: c <= 9'b101101100;
				8'b1110101: c <= 9'b101110000;
				8'b1111101: c <= 9'b111110101;
				8'b101001: c <= 9'b111000010;
				8'b1010010: c <= 9'b100111000;
				8'b1011000: c <= 9'b110000101;
				8'b101110: c <= 9'b11010111;
				8'b1000001: c <= 9'b1000000;
				default: c <= 9'b0;
			endcase
			9'b100110110 : case(di)
				8'b1000011: c <= 9'b1100110;
				8'b101000: c <= 9'b1010010;
				8'b111010: c <= 9'b111111111;
				8'b110110: c <= 9'b111110000;
				8'b1100100: c <= 9'b1001;
				8'b1000000: c <= 9'b11101100;
				8'b1110110: c <= 9'b11101111;
				8'b100101: c <= 9'b111011111;
				8'b101111: c <= 9'b10111010;
				8'b100110: c <= 9'b11001011;
				8'b1100011: c <= 9'b10001100;
				8'b1001000: c <= 9'b111000100;
				8'b111000: c <= 9'b111111;
				8'b110001: c <= 9'b1001010;
				8'b1010111: c <= 9'b10100101;
				8'b1001110: c <= 9'b101010010;
				8'b1101010: c <= 9'b101110100;
				8'b1001001: c <= 9'b100011100;
				8'b1100000: c <= 9'b110001101;
				8'b110111: c <= 9'b111000000;
				8'b1011101: c <= 9'b110101;
				8'b1011011: c <= 9'b110110110;
				8'b111001: c <= 9'b11100010;
				8'b1001010: c <= 9'b11000110;
				8'b110011: c <= 9'b1011100;
				8'b1101100: c <= 9'b11001;
				8'b1110111: c <= 9'b10100111;
				8'b101011: c <= 9'b10000111;
				8'b1101011: c <= 9'b110001011;
				8'b111100: c <= 9'b1011000;
				8'b1000111: c <= 9'b10110111;
				8'b1011111: c <= 9'b111000011;
				8'b1110100: c <= 9'b100010111;
				8'b101101: c <= 9'b11011;
				8'b1010011: c <= 9'b100110010;
				8'b1100001: c <= 9'b111000011;
				8'b110101: c <= 9'b100010000;
				8'b1000100: c <= 9'b111;
				8'b1010001: c <= 9'b10111101;
				8'b1010100: c <= 9'b110111010;
				8'b1100110: c <= 9'b111101111;
				8'b101010: c <= 9'b110110110;
				8'b1011110: c <= 9'b100010000;
				8'b1100111: c <= 9'b1110;
				8'b1011010: c <= 9'b10111011;
				8'b1000010: c <= 9'b110100;
				8'b111101: c <= 9'b111101;
				8'b110000: c <= 9'b100100101;
				8'b111110: c <= 9'b101000001;
				8'b1100010: c <= 9'b110101011;
				8'b1110000: c <= 9'b101101101;
				8'b1101001: c <= 9'b101101101;
				8'b1110011: c <= 9'b101101100;
				8'b1001100: c <= 9'b10010011;
				8'b100001: c <= 9'b11011000;
				8'b1000110: c <= 9'b101000100;
				8'b1110010: c <= 9'b111000010;
				8'b1010000: c <= 9'b100111110;
				8'b1111010: c <= 9'b101101011;
				8'b1010101: c <= 9'b1101101;
				8'b111011: c <= 9'b100100;
				8'b1001101: c <= 9'b101011101;
				8'b111111: c <= 9'b110011000;
				8'b1101110: c <= 9'b10101001;
				8'b1111011: c <= 9'b111001110;
				8'b1001011: c <= 9'b11101100;
				8'b1101111: c <= 9'b100011101;
				8'b1101000: c <= 9'b10000111;
				8'b101100: c <= 9'b10011000;
				8'b100100: c <= 9'b111010110;
				8'b1111000: c <= 9'b10111111;
				8'b1000101: c <= 9'b100001111;
				8'b1011001: c <= 9'b101011;
				8'b110100: c <= 9'b110110100;
				8'b1111001: c <= 9'b111;
				8'b1110001: c <= 9'b101111001;
				8'b1001111: c <= 9'b10001111;
				8'b1100101: c <= 9'b100001100;
				8'b1111110: c <= 9'b1110;
				8'b1111100: c <= 9'b11100100;
				8'b1010110: c <= 9'b10000110;
				8'b110010: c <= 9'b11100110;
				8'b1101101: c <= 9'b10011001;
				8'b100011: c <= 9'b100110;
				8'b1110101: c <= 9'b101110111;
				8'b1111101: c <= 9'b110110100;
				8'b101001: c <= 9'b101110000;
				8'b1010010: c <= 9'b101001100;
				8'b1011000: c <= 9'b101011010;
				8'b101110: c <= 9'b1010000;
				8'b1000001: c <= 9'b11100010;
				default: c <= 9'b0;
			endcase
			9'b1101000 : case(di)
				8'b1000011: c <= 9'b11010101;
				8'b101000: c <= 9'b1110;
				8'b111010: c <= 9'b101101000;
				8'b110110: c <= 9'b11101101;
				8'b1100100: c <= 9'b100010001;
				8'b1000000: c <= 9'b110011111;
				8'b1110110: c <= 9'b11100101;
				8'b100101: c <= 9'b101111110;
				8'b101111: c <= 9'b11100110;
				8'b100110: c <= 9'b110011;
				8'b1100011: c <= 9'b100101101;
				8'b1001000: c <= 9'b100110111;
				8'b111000: c <= 9'b101001010;
				8'b110001: c <= 9'b111011110;
				8'b1010111: c <= 9'b10011000;
				8'b1001110: c <= 9'b110110;
				8'b1101010: c <= 9'b100110110;
				8'b1001001: c <= 9'b101001000;
				8'b1100000: c <= 9'b10;
				8'b110111: c <= 9'b110110010;
				8'b1011101: c <= 9'b101001010;
				8'b1011011: c <= 9'b10111010;
				8'b111001: c <= 9'b10111;
				8'b1001010: c <= 9'b1110;
				8'b110011: c <= 9'b110000111;
				8'b1101100: c <= 9'b1001000;
				8'b1110111: c <= 9'b1110101;
				8'b101011: c <= 9'b100001101;
				8'b1101011: c <= 9'b11101000;
				8'b111100: c <= 9'b10000001;
				8'b1000111: c <= 9'b10110;
				8'b1011111: c <= 9'b101110010;
				8'b1110100: c <= 9'b101010011;
				8'b101101: c <= 9'b110001110;
				8'b1010011: c <= 9'b101001010;
				8'b1100001: c <= 9'b10100111;
				8'b110101: c <= 9'b101101010;
				8'b1000100: c <= 9'b101110011;
				8'b1010001: c <= 9'b101010;
				8'b1010100: c <= 9'b111100000;
				8'b1100110: c <= 9'b111010100;
				8'b101010: c <= 9'b110110111;
				8'b1011110: c <= 9'b11100100;
				8'b1100111: c <= 9'b11011011;
				8'b1011010: c <= 9'b110010111;
				8'b1000010: c <= 9'b11000010;
				8'b111101: c <= 9'b101100100;
				8'b110000: c <= 9'b110111110;
				8'b111110: c <= 9'b11000011;
				8'b1100010: c <= 9'b11110110;
				8'b1110000: c <= 9'b11101000;
				8'b1101001: c <= 9'b111111000;
				8'b1110011: c <= 9'b111001000;
				8'b1001100: c <= 9'b11011011;
				8'b100001: c <= 9'b101110101;
				8'b1000110: c <= 9'b1100010;
				8'b1110010: c <= 9'b111010010;
				8'b1010000: c <= 9'b100100011;
				8'b1111010: c <= 9'b10101010;
				8'b1010101: c <= 9'b10101;
				8'b111011: c <= 9'b11001001;
				8'b1001101: c <= 9'b1011000;
				8'b111111: c <= 9'b1011111;
				8'b1101110: c <= 9'b110000;
				8'b1111011: c <= 9'b110100000;
				8'b1001011: c <= 9'b1110001;
				8'b1101111: c <= 9'b1001;
				8'b1101000: c <= 9'b1100011;
				8'b101100: c <= 9'b10110011;
				8'b100100: c <= 9'b110100010;
				8'b1111000: c <= 9'b100111100;
				8'b1000101: c <= 9'b110010;
				8'b1011001: c <= 9'b11011100;
				8'b110100: c <= 9'b111011111;
				8'b1111001: c <= 9'b110100100;
				8'b1110001: c <= 9'b1110101;
				8'b1001111: c <= 9'b10111110;
				8'b1100101: c <= 9'b110110101;
				8'b1111110: c <= 9'b11001001;
				8'b1111100: c <= 9'b100110110;
				8'b1010110: c <= 9'b100001111;
				8'b110010: c <= 9'b10101100;
				8'b1101101: c <= 9'b101011111;
				8'b100011: c <= 9'b100011011;
				8'b1110101: c <= 9'b1111010;
				8'b1111101: c <= 9'b100010111;
				8'b101001: c <= 9'b101001110;
				8'b1010010: c <= 9'b1111;
				8'b1011000: c <= 9'b111011010;
				8'b101110: c <= 9'b101110110;
				8'b1000001: c <= 9'b10111;
				default: c <= 9'b0;
			endcase
			9'b110001100 : case(di)
				8'b1000011: c <= 9'b1001010;
				8'b101000: c <= 9'b111011011;
				8'b111010: c <= 9'b100011010;
				8'b110110: c <= 9'b11001111;
				8'b1100100: c <= 9'b10010101;
				8'b1000000: c <= 9'b1000100;
				8'b1110110: c <= 9'b11011000;
				8'b100101: c <= 9'b11010111;
				8'b101111: c <= 9'b11010111;
				8'b100110: c <= 9'b100110110;
				8'b1100011: c <= 9'b11100100;
				8'b1001000: c <= 9'b11001000;
				8'b111000: c <= 9'b10101100;
				8'b110001: c <= 9'b110101111;
				8'b1010111: c <= 9'b100001101;
				8'b1001110: c <= 9'b11100010;
				8'b1101010: c <= 9'b101000111;
				8'b1001001: c <= 9'b11000011;
				8'b1100000: c <= 9'b110001000;
				8'b110111: c <= 9'b100000011;
				8'b1011101: c <= 9'b1101100;
				8'b1011011: c <= 9'b10111000;
				8'b111001: c <= 9'b111101101;
				8'b1001010: c <= 9'b100100000;
				8'b110011: c <= 9'b100011000;
				8'b1101100: c <= 9'b10011011;
				8'b1110111: c <= 9'b1110011;
				8'b101011: c <= 9'b101110110;
				8'b1101011: c <= 9'b111001011;
				8'b111100: c <= 9'b101100101;
				8'b1000111: c <= 9'b10010;
				8'b1011111: c <= 9'b110;
				8'b1110100: c <= 9'b11100110;
				8'b101101: c <= 9'b111111110;
				8'b1010011: c <= 9'b100001101;
				8'b1100001: c <= 9'b111000000;
				8'b110101: c <= 9'b11110010;
				8'b1000100: c <= 9'b10100100;
				8'b1010001: c <= 9'b111011100;
				8'b1010100: c <= 9'b10001011;
				8'b1100110: c <= 9'b100011001;
				8'b101010: c <= 9'b110010110;
				8'b1011110: c <= 9'b101100101;
				8'b1100111: c <= 9'b110001101;
				8'b1011010: c <= 9'b111000110;
				8'b1000010: c <= 9'b100001010;
				8'b111101: c <= 9'b1111101;
				8'b110000: c <= 9'b100010110;
				8'b111110: c <= 9'b10111010;
				8'b1100010: c <= 9'b1001001;
				8'b1110000: c <= 9'b100001;
				8'b1101001: c <= 9'b10010100;
				8'b1110011: c <= 9'b100101111;
				8'b1001100: c <= 9'b111001001;
				8'b100001: c <= 9'b101011;
				8'b1000110: c <= 9'b100101011;
				8'b1110010: c <= 9'b111000111;
				8'b1010000: c <= 9'b100001100;
				8'b1111010: c <= 9'b100001111;
				8'b1010101: c <= 9'b10111010;
				8'b111011: c <= 9'b111011011;
				8'b1001101: c <= 9'b100100000;
				8'b111111: c <= 9'b1100111;
				8'b1101110: c <= 9'b111100110;
				8'b1111011: c <= 9'b11011101;
				8'b1001011: c <= 9'b111001110;
				8'b1101111: c <= 9'b1010010;
				8'b1101000: c <= 9'b1010101;
				8'b101100: c <= 9'b1010000;
				8'b100100: c <= 9'b111000010;
				8'b1111000: c <= 9'b10111011;
				8'b1000101: c <= 9'b111000111;
				8'b1011001: c <= 9'b110001000;
				8'b110100: c <= 9'b100101000;
				8'b1111001: c <= 9'b110000011;
				8'b1110001: c <= 9'b10100010;
				8'b1001111: c <= 9'b111100001;
				8'b1100101: c <= 9'b111010110;
				8'b1111110: c <= 9'b111111011;
				8'b1111100: c <= 9'b111011111;
				8'b1010110: c <= 9'b111000101;
				8'b110010: c <= 9'b101000100;
				8'b1101101: c <= 9'b100001001;
				8'b100011: c <= 9'b101111111;
				8'b1110101: c <= 9'b11100000;
				8'b1111101: c <= 9'b110100;
				8'b101001: c <= 9'b111001;
				8'b1010010: c <= 9'b110010001;
				8'b1011000: c <= 9'b100010000;
				8'b101110: c <= 9'b110011010;
				8'b1000001: c <= 9'b1100000;
				default: c <= 9'b0;
			endcase
			9'b11000000 : case(di)
				8'b1000011: c <= 9'b100111101;
				8'b101000: c <= 9'b100001101;
				8'b111010: c <= 9'b10100010;
				8'b110110: c <= 9'b10001110;
				8'b1100100: c <= 9'b10111001;
				8'b1000000: c <= 9'b11110010;
				8'b1110110: c <= 9'b10000;
				8'b100101: c <= 9'b110000;
				8'b101111: c <= 9'b110001100;
				8'b100110: c <= 9'b100010101;
				8'b1100011: c <= 9'b100100010;
				8'b1001000: c <= 9'b100101111;
				8'b111000: c <= 9'b111111011;
				8'b110001: c <= 9'b100000111;
				8'b1010111: c <= 9'b110010110;
				8'b1001110: c <= 9'b100001101;
				8'b1101010: c <= 9'b101110100;
				8'b1001001: c <= 9'b110010100;
				8'b1100000: c <= 9'b111011010;
				8'b110111: c <= 9'b10100;
				8'b1011101: c <= 9'b11011100;
				8'b1011011: c <= 9'b100110110;
				8'b111001: c <= 9'b1101110;
				8'b1001010: c <= 9'b101010000;
				8'b110011: c <= 9'b101110;
				8'b1101100: c <= 9'b1001;
				8'b1110111: c <= 9'b111000100;
				8'b101011: c <= 9'b111011110;
				8'b1101011: c <= 9'b110110100;
				8'b111100: c <= 9'b10001101;
				8'b1000111: c <= 9'b11010101;
				8'b1011111: c <= 9'b111001110;
				8'b1110100: c <= 9'b101100011;
				8'b101101: c <= 9'b100000100;
				8'b1010011: c <= 9'b1001;
				8'b1100001: c <= 9'b101011;
				8'b110101: c <= 9'b101101111;
				8'b1000100: c <= 9'b110011;
				8'b1010001: c <= 9'b101100011;
				8'b1010100: c <= 9'b1100100;
				8'b1100110: c <= 9'b100100110;
				8'b101010: c <= 9'b1011000;
				8'b1011110: c <= 9'b11111101;
				8'b1100111: c <= 9'b10100110;
				8'b1011010: c <= 9'b100011011;
				8'b1000010: c <= 9'b10101001;
				8'b111101: c <= 9'b110001010;
				8'b110000: c <= 9'b110101010;
				8'b111110: c <= 9'b101111111;
				8'b1100010: c <= 9'b100001111;
				8'b1110000: c <= 9'b1101;
				8'b1101001: c <= 9'b1100001;
				8'b1110011: c <= 9'b111000010;
				8'b1001100: c <= 9'b110111111;
				8'b100001: c <= 9'b10111;
				8'b1000110: c <= 9'b111001;
				8'b1110010: c <= 9'b11110111;
				8'b1010000: c <= 9'b100111111;
				8'b1111010: c <= 9'b1110011;
				8'b1010101: c <= 9'b10010000;
				8'b111011: c <= 9'b10101001;
				8'b1001101: c <= 9'b1000001;
				8'b111111: c <= 9'b110000011;
				8'b1101110: c <= 9'b100100001;
				8'b1111011: c <= 9'b1010011;
				8'b1001011: c <= 9'b110011010;
				8'b1101111: c <= 9'b100001111;
				8'b1101000: c <= 9'b111000111;
				8'b101100: c <= 9'b10011011;
				8'b100100: c <= 9'b100001111;
				8'b1111000: c <= 9'b101010101;
				8'b1000101: c <= 9'b1110010;
				8'b1011001: c <= 9'b100101000;
				8'b110100: c <= 9'b101010111;
				8'b1111001: c <= 9'b101011011;
				8'b1110001: c <= 9'b110110;
				8'b1001111: c <= 9'b1101101;
				8'b1100101: c <= 9'b100101110;
				8'b1111110: c <= 9'b10010101;
				8'b1111100: c <= 9'b110001011;
				8'b1010110: c <= 9'b1111010;
				8'b110010: c <= 9'b101;
				8'b1101101: c <= 9'b11011101;
				8'b100011: c <= 9'b111101100;
				8'b1110101: c <= 9'b101010001;
				8'b1111101: c <= 9'b111100110;
				8'b101001: c <= 9'b10111111;
				8'b1010010: c <= 9'b1101101;
				8'b1011000: c <= 9'b1111101;
				8'b101110: c <= 9'b111010100;
				8'b1000001: c <= 9'b101001010;
				default: c <= 9'b0;
			endcase
			9'b111011001 : case(di)
				8'b1000011: c <= 9'b111111;
				8'b101000: c <= 9'b100;
				8'b111010: c <= 9'b100101101;
				8'b110110: c <= 9'b101011101;
				8'b1100100: c <= 9'b11100110;
				8'b1000000: c <= 9'b100001101;
				8'b1110110: c <= 9'b1011010;
				8'b100101: c <= 9'b1101100;
				8'b101111: c <= 9'b10000101;
				8'b100110: c <= 9'b10111010;
				8'b1100011: c <= 9'b10010;
				8'b1001000: c <= 9'b110100101;
				8'b111000: c <= 9'b100101101;
				8'b110001: c <= 9'b1101000;
				8'b1010111: c <= 9'b110101011;
				8'b1001110: c <= 9'b1111100;
				8'b1101010: c <= 9'b110100010;
				8'b1001001: c <= 9'b101111110;
				8'b1100000: c <= 9'b11111011;
				8'b110111: c <= 9'b100110;
				8'b1011101: c <= 9'b100110111;
				8'b1011011: c <= 9'b111110101;
				8'b111001: c <= 9'b110011100;
				8'b1001010: c <= 9'b100000011;
				8'b110011: c <= 9'b11101000;
				8'b1101100: c <= 9'b11011101;
				8'b1110111: c <= 9'b111101000;
				8'b101011: c <= 9'b111011101;
				8'b1101011: c <= 9'b1101000;
				8'b111100: c <= 9'b101110001;
				8'b1000111: c <= 9'b10001001;
				8'b1011111: c <= 9'b100101001;
				8'b1110100: c <= 9'b110001111;
				8'b101101: c <= 9'b101010000;
				8'b1010011: c <= 9'b11000;
				8'b1100001: c <= 9'b111001001;
				8'b110101: c <= 9'b1001101;
				8'b1000100: c <= 9'b100110010;
				8'b1010001: c <= 9'b1111100;
				8'b1010100: c <= 9'b10010001;
				8'b1100110: c <= 9'b10010;
				8'b101010: c <= 9'b100011111;
				8'b1011110: c <= 9'b100101;
				8'b1100111: c <= 9'b10011111;
				8'b1011010: c <= 9'b110111110;
				8'b1000010: c <= 9'b100110100;
				8'b111101: c <= 9'b100110000;
				8'b110000: c <= 9'b111001001;
				8'b111110: c <= 9'b10001001;
				8'b1100010: c <= 9'b111010110;
				8'b1110000: c <= 9'b110000;
				8'b1101001: c <= 9'b100110011;
				8'b1110011: c <= 9'b101110110;
				8'b1001100: c <= 9'b111000000;
				8'b100001: c <= 9'b1110;
				8'b1000110: c <= 9'b101010000;
				8'b1110010: c <= 9'b110100001;
				8'b1010000: c <= 9'b100001011;
				8'b1111010: c <= 9'b111010100;
				8'b1010101: c <= 9'b10010001;
				8'b111011: c <= 9'b1001111;
				8'b1001101: c <= 9'b1111;
				8'b111111: c <= 9'b100001100;
				8'b1101110: c <= 9'b1;
				8'b1111011: c <= 9'b110001010;
				8'b1001011: c <= 9'b1010001;
				8'b1101111: c <= 9'b110100111;
				8'b1101000: c <= 9'b101000100;
				8'b101100: c <= 9'b101011010;
				8'b100100: c <= 9'b101011000;
				8'b1111000: c <= 9'b100100;
				8'b1000101: c <= 9'b111101111;
				8'b1011001: c <= 9'b100110100;
				8'b110100: c <= 9'b11011101;
				8'b1111001: c <= 9'b1101101;
				8'b1110001: c <= 9'b11010111;
				8'b1001111: c <= 9'b101000;
				8'b1100101: c <= 9'b100010011;
				8'b1111110: c <= 9'b10;
				8'b1111100: c <= 9'b111011101;
				8'b1010110: c <= 9'b1101000;
				8'b110010: c <= 9'b100000111;
				8'b1101101: c <= 9'b101100001;
				8'b100011: c <= 9'b100111000;
				8'b1110101: c <= 9'b10111111;
				8'b1111101: c <= 9'b101101000;
				8'b101001: c <= 9'b11100010;
				8'b1010010: c <= 9'b1100101;
				8'b1011000: c <= 9'b1110100;
				8'b101110: c <= 9'b11001011;
				8'b1000001: c <= 9'b100001;
				default: c <= 9'b0;
			endcase
			9'b110001011 : case(di)
				8'b1000011: c <= 9'b111010010;
				8'b101000: c <= 9'b1000101;
				8'b111010: c <= 9'b11101111;
				8'b110110: c <= 9'b100100000;
				8'b1100100: c <= 9'b101101010;
				8'b1000000: c <= 9'b1100111;
				8'b1110110: c <= 9'b11000000;
				8'b100101: c <= 9'b110111011;
				8'b101111: c <= 9'b100111001;
				8'b100110: c <= 9'b11110101;
				8'b1100011: c <= 9'b100011100;
				8'b1001000: c <= 9'b100011101;
				8'b111000: c <= 9'b11101000;
				8'b110001: c <= 9'b1100101;
				8'b1010111: c <= 9'b110111011;
				8'b1001110: c <= 9'b110100111;
				8'b1101010: c <= 9'b110000000;
				8'b1001001: c <= 9'b101000111;
				8'b1100000: c <= 9'b11;
				8'b110111: c <= 9'b111111;
				8'b1011101: c <= 9'b11010;
				8'b1011011: c <= 9'b111001100;
				8'b111001: c <= 9'b110001001;
				8'b1001010: c <= 9'b1000011;
				8'b110011: c <= 9'b11100100;
				8'b1101100: c <= 9'b100110110;
				8'b1110111: c <= 9'b1000100;
				8'b101011: c <= 9'b10000001;
				8'b1101011: c <= 9'b110110110;
				8'b111100: c <= 9'b101011110;
				8'b1000111: c <= 9'b11011001;
				8'b1011111: c <= 9'b111100001;
				8'b1110100: c <= 9'b10011011;
				8'b101101: c <= 9'b111111;
				8'b1010011: c <= 9'b1101001;
				8'b1100001: c <= 9'b110101010;
				8'b110101: c <= 9'b100101010;
				8'b1000100: c <= 9'b110011101;
				8'b1010001: c <= 9'b1001110;
				8'b1010100: c <= 9'b101110111;
				8'b1100110: c <= 9'b11000000;
				8'b101010: c <= 9'b111011101;
				8'b1011110: c <= 9'b101111010;
				8'b1100111: c <= 9'b11100111;
				8'b1011010: c <= 9'b101011011;
				8'b1000010: c <= 9'b1000011;
				8'b111101: c <= 9'b1100001;
				8'b110000: c <= 9'b11101011;
				8'b111110: c <= 9'b11001100;
				8'b1100010: c <= 9'b1001101;
				8'b1110000: c <= 9'b100001100;
				8'b1101001: c <= 9'b110100110;
				8'b1110011: c <= 9'b101000100;
				8'b1001100: c <= 9'b101110;
				8'b100001: c <= 9'b101111111;
				8'b1000110: c <= 9'b100011010;
				8'b1110010: c <= 9'b111101010;
				8'b1010000: c <= 9'b11100;
				8'b1111010: c <= 9'b111110000;
				8'b1010101: c <= 9'b111011111;
				8'b111011: c <= 9'b100010011;
				8'b1001101: c <= 9'b111100010;
				8'b111111: c <= 9'b100110000;
				8'b1101110: c <= 9'b101100000;
				8'b1111011: c <= 9'b111100111;
				8'b1001011: c <= 9'b101110001;
				8'b1101111: c <= 9'b111111010;
				8'b1101000: c <= 9'b100101110;
				8'b101100: c <= 9'b110011;
				8'b100100: c <= 9'b111100;
				8'b1111000: c <= 9'b10010000;
				8'b1000101: c <= 9'b10000110;
				8'b1011001: c <= 9'b10110;
				8'b110100: c <= 9'b10101100;
				8'b1111001: c <= 9'b10101111;
				8'b1110001: c <= 9'b11010001;
				8'b1001111: c <= 9'b101000001;
				8'b1100101: c <= 9'b110100100;
				8'b1111110: c <= 9'b101011011;
				8'b1111100: c <= 9'b101010;
				8'b1010110: c <= 9'b101000011;
				8'b110010: c <= 9'b101001111;
				8'b1101101: c <= 9'b10101100;
				8'b100011: c <= 9'b110111;
				8'b1110101: c <= 9'b1001000;
				8'b1111101: c <= 9'b10110010;
				8'b101001: c <= 9'b10000110;
				8'b1010010: c <= 9'b11100011;
				8'b1011000: c <= 9'b110110111;
				8'b101110: c <= 9'b11000111;
				8'b1000001: c <= 9'b100001011;
				default: c <= 9'b0;
			endcase
			9'b101101010 : case(di)
				8'b1000011: c <= 9'b111101111;
				8'b101000: c <= 9'b10011011;
				8'b111010: c <= 9'b10110111;
				8'b110110: c <= 9'b10111000;
				8'b1100100: c <= 9'b11;
				8'b1000000: c <= 9'b1101100;
				8'b1110110: c <= 9'b111000101;
				8'b100101: c <= 9'b101101100;
				8'b101111: c <= 9'b100110010;
				8'b100110: c <= 9'b11100110;
				8'b1100011: c <= 9'b110110010;
				8'b1001000: c <= 9'b110001;
				8'b111000: c <= 9'b110001101;
				8'b110001: c <= 9'b101110101;
				8'b1010111: c <= 9'b101010011;
				8'b1001110: c <= 9'b1001101;
				8'b1101010: c <= 9'b100010100;
				8'b1001001: c <= 9'b10000101;
				8'b1100000: c <= 9'b10001101;
				8'b110111: c <= 9'b101001011;
				8'b1011101: c <= 9'b111011111;
				8'b1011011: c <= 9'b111001111;
				8'b111001: c <= 9'b1110111;
				8'b1001010: c <= 9'b111010110;
				8'b110011: c <= 9'b10010110;
				8'b1101100: c <= 9'b10000010;
				8'b1110111: c <= 9'b1000110;
				8'b101011: c <= 9'b101010000;
				8'b1101011: c <= 9'b100110;
				8'b111100: c <= 9'b11101;
				8'b1000111: c <= 9'b111110110;
				8'b1011111: c <= 9'b111000111;
				8'b1110100: c <= 9'b111000110;
				8'b101101: c <= 9'b1001000;
				8'b1010011: c <= 9'b11000000;
				8'b1100001: c <= 9'b100001100;
				8'b110101: c <= 9'b111011110;
				8'b1000100: c <= 9'b101100011;
				8'b1010001: c <= 9'b100111100;
				8'b1010100: c <= 9'b1010101;
				8'b1100110: c <= 9'b10000110;
				8'b101010: c <= 9'b11110110;
				8'b1011110: c <= 9'b1100111;
				8'b1100111: c <= 9'b10011;
				8'b1011010: c <= 9'b1110101;
				8'b1000010: c <= 9'b110111011;
				8'b111101: c <= 9'b11101011;
				8'b110000: c <= 9'b10100;
				8'b111110: c <= 9'b111011111;
				8'b1100010: c <= 9'b1001;
				8'b1110000: c <= 9'b110111011;
				8'b1101001: c <= 9'b101000;
				8'b1110011: c <= 9'b110100101;
				8'b1001100: c <= 9'b11110100;
				8'b100001: c <= 9'b11100;
				8'b1000110: c <= 9'b110110100;
				8'b1110010: c <= 9'b11011;
				8'b1010000: c <= 9'b10000111;
				8'b1111010: c <= 9'b10111101;
				8'b1010101: c <= 9'b111100010;
				8'b111011: c <= 9'b101110011;
				8'b1001101: c <= 9'b11001;
				8'b111111: c <= 9'b100010110;
				8'b1101110: c <= 9'b101010001;
				8'b1111011: c <= 9'b10111000;
				8'b1001011: c <= 9'b11111;
				8'b1101111: c <= 9'b111010000;
				8'b1101000: c <= 9'b111110101;
				8'b101100: c <= 9'b11101101;
				8'b100100: c <= 9'b11110110;
				8'b1111000: c <= 9'b111010110;
				8'b1000101: c <= 9'b10011101;
				8'b1011001: c <= 9'b10101011;
				8'b110100: c <= 9'b100010011;
				8'b1111001: c <= 9'b111001101;
				8'b1110001: c <= 9'b111101010;
				8'b1001111: c <= 9'b11000001;
				8'b1100101: c <= 9'b11101001;
				8'b1111110: c <= 9'b111111011;
				8'b1111100: c <= 9'b100100101;
				8'b1010110: c <= 9'b1011000;
				8'b110010: c <= 9'b100010010;
				8'b1101101: c <= 9'b1101;
				8'b100011: c <= 9'b110011001;
				8'b1110101: c <= 9'b10101011;
				8'b1111101: c <= 9'b110001110;
				8'b101001: c <= 9'b101111010;
				8'b1010010: c <= 9'b101010011;
				8'b1011000: c <= 9'b100101110;
				8'b101110: c <= 9'b101011011;
				8'b1000001: c <= 9'b11000111;
				default: c <= 9'b0;
			endcase
			9'b111001011 : case(di)
				8'b1000011: c <= 9'b10011001;
				8'b101000: c <= 9'b10;
				8'b111010: c <= 9'b110010101;
				8'b110110: c <= 9'b101000;
				8'b1100100: c <= 9'b11110101;
				8'b1000000: c <= 9'b100110010;
				8'b1110110: c <= 9'b101100100;
				8'b100101: c <= 9'b1110011;
				8'b101111: c <= 9'b111010;
				8'b100110: c <= 9'b110100;
				8'b1100011: c <= 9'b111001;
				8'b1001000: c <= 9'b110110010;
				8'b111000: c <= 9'b101100001;
				8'b110001: c <= 9'b101010110;
				8'b1010111: c <= 9'b11111011;
				8'b1001110: c <= 9'b111111011;
				8'b1101010: c <= 9'b100000000;
				8'b1001001: c <= 9'b100100011;
				8'b1100000: c <= 9'b101100100;
				8'b110111: c <= 9'b100000101;
				8'b1011101: c <= 9'b11110000;
				8'b1011011: c <= 9'b100010101;
				8'b111001: c <= 9'b10111001;
				8'b1001010: c <= 9'b10111001;
				8'b110011: c <= 9'b100010000;
				8'b1101100: c <= 9'b101111110;
				8'b1110111: c <= 9'b1001111;
				8'b101011: c <= 9'b10101101;
				8'b1101011: c <= 9'b10001110;
				8'b111100: c <= 9'b11111001;
				8'b1000111: c <= 9'b111100001;
				8'b1011111: c <= 9'b100001110;
				8'b1110100: c <= 9'b111001010;
				8'b101101: c <= 9'b110001111;
				8'b1010011: c <= 9'b110011000;
				8'b1100001: c <= 9'b101111110;
				8'b110101: c <= 9'b10100110;
				8'b1000100: c <= 9'b10100010;
				8'b1010001: c <= 9'b101110000;
				8'b1010100: c <= 9'b110100011;
				8'b1100110: c <= 9'b101010000;
				8'b101010: c <= 9'b100011100;
				8'b1011110: c <= 9'b10111010;
				8'b1100111: c <= 9'b110101111;
				8'b1011010: c <= 9'b1001110;
				8'b1000010: c <= 9'b111110110;
				8'b111101: c <= 9'b111000101;
				8'b110000: c <= 9'b1000000;
				8'b111110: c <= 9'b11011001;
				8'b1100010: c <= 9'b1011001;
				8'b1110000: c <= 9'b1100111;
				8'b1101001: c <= 9'b101000010;
				8'b1110011: c <= 9'b111100100;
				8'b1001100: c <= 9'b1001000;
				8'b100001: c <= 9'b100110111;
				8'b1000110: c <= 9'b1001000;
				8'b1110010: c <= 9'b11101101;
				8'b1010000: c <= 9'b100010000;
				8'b1111010: c <= 9'b1110011;
				8'b1010101: c <= 9'b1001101;
				8'b111011: c <= 9'b100100111;
				8'b1001101: c <= 9'b11110110;
				8'b111111: c <= 9'b11101000;
				8'b1101110: c <= 9'b1111011;
				8'b1111011: c <= 9'b110100010;
				8'b1001011: c <= 9'b11010011;
				8'b1101111: c <= 9'b1111011;
				8'b1101000: c <= 9'b100001010;
				8'b101100: c <= 9'b11100011;
				8'b100100: c <= 9'b100010101;
				8'b1111000: c <= 9'b10000;
				8'b1000101: c <= 9'b1;
				8'b1011001: c <= 9'b110111100;
				8'b110100: c <= 9'b110001010;
				8'b1111001: c <= 9'b110000011;
				8'b1110001: c <= 9'b110111100;
				8'b1001111: c <= 9'b100101110;
				8'b1100101: c <= 9'b100111110;
				8'b1111110: c <= 9'b10000111;
				8'b1111100: c <= 9'b100100111;
				8'b1010110: c <= 9'b101010011;
				8'b110010: c <= 9'b111110101;
				8'b1101101: c <= 9'b111111110;
				8'b100011: c <= 9'b10100110;
				8'b1110101: c <= 9'b11110;
				8'b1111101: c <= 9'b11111101;
				8'b101001: c <= 9'b111011;
				8'b1010010: c <= 9'b101110000;
				8'b1011000: c <= 9'b110000111;
				8'b101110: c <= 9'b10111111;
				8'b1000001: c <= 9'b11000001;
				default: c <= 9'b0;
			endcase
			9'b111100101 : case(di)
				8'b1000011: c <= 9'b11111011;
				8'b101000: c <= 9'b10001101;
				8'b111010: c <= 9'b110010101;
				8'b110110: c <= 9'b100110101;
				8'b1100100: c <= 9'b1011110;
				8'b1000000: c <= 9'b11010011;
				8'b1110110: c <= 9'b10010011;
				8'b100101: c <= 9'b101001011;
				8'b101111: c <= 9'b111101;
				8'b100110: c <= 9'b101000011;
				8'b1100011: c <= 9'b111000010;
				8'b1001000: c <= 9'b10001100;
				8'b111000: c <= 9'b111001111;
				8'b110001: c <= 9'b110011000;
				8'b1010111: c <= 9'b10110010;
				8'b1001110: c <= 9'b10100110;
				8'b1101010: c <= 9'b11001100;
				8'b1001001: c <= 9'b10111101;
				8'b1100000: c <= 9'b111000101;
				8'b110111: c <= 9'b100001011;
				8'b1011101: c <= 9'b101110110;
				8'b1011011: c <= 9'b110001011;
				8'b111001: c <= 9'b110001100;
				8'b1001010: c <= 9'b1001000;
				8'b110011: c <= 9'b110101001;
				8'b1101100: c <= 9'b110100000;
				8'b1110111: c <= 9'b11100001;
				8'b101011: c <= 9'b101010000;
				8'b1101011: c <= 9'b11010010;
				8'b111100: c <= 9'b111110101;
				8'b1000111: c <= 9'b1100;
				8'b1011111: c <= 9'b10001100;
				8'b1110100: c <= 9'b100100110;
				8'b101101: c <= 9'b10000011;
				8'b1010011: c <= 9'b1000010;
				8'b1100001: c <= 9'b110000101;
				8'b110101: c <= 9'b100011010;
				8'b1000100: c <= 9'b10;
				8'b1010001: c <= 9'b110001;
				8'b1010100: c <= 9'b1001010;
				8'b1100110: c <= 9'b11101000;
				8'b101010: c <= 9'b101110111;
				8'b1011110: c <= 9'b10100100;
				8'b1100111: c <= 9'b111001111;
				8'b1011010: c <= 9'b1001101;
				8'b1000010: c <= 9'b100000111;
				8'b111101: c <= 9'b101001011;
				8'b110000: c <= 9'b110111010;
				8'b111110: c <= 9'b1011011;
				8'b1100010: c <= 9'b100001100;
				8'b1110000: c <= 9'b100100010;
				8'b1101001: c <= 9'b110100;
				8'b1110011: c <= 9'b100010;
				8'b1001100: c <= 9'b110001010;
				8'b100001: c <= 9'b100000010;
				8'b1000110: c <= 9'b111110011;
				8'b1110010: c <= 9'b110011010;
				8'b1010000: c <= 9'b101;
				8'b1111010: c <= 9'b11001011;
				8'b1010101: c <= 9'b11101111;
				8'b111011: c <= 9'b11101001;
				8'b1001101: c <= 9'b1111001;
				8'b111111: c <= 9'b11011101;
				8'b1101110: c <= 9'b100;
				8'b1111011: c <= 9'b10100110;
				8'b1001011: c <= 9'b10011001;
				8'b1101111: c <= 9'b101011011;
				8'b1101000: c <= 9'b10101101;
				8'b101100: c <= 9'b100100011;
				8'b100100: c <= 9'b10101011;
				8'b1111000: c <= 9'b100001110;
				8'b1000101: c <= 9'b1001011;
				8'b1011001: c <= 9'b1000101;
				8'b110100: c <= 9'b101001;
				8'b1111001: c <= 9'b10101111;
				8'b1110001: c <= 9'b111001111;
				8'b1001111: c <= 9'b111101111;
				8'b1100101: c <= 9'b100011010;
				8'b1111110: c <= 9'b10010;
				8'b1111100: c <= 9'b1000000;
				8'b1010110: c <= 9'b101000100;
				8'b110010: c <= 9'b10000001;
				8'b1101101: c <= 9'b111100101;
				8'b100011: c <= 9'b100001;
				8'b1110101: c <= 9'b101100010;
				8'b1111101: c <= 9'b111011101;
				8'b101001: c <= 9'b1111000;
				8'b1010010: c <= 9'b1000100;
				8'b1011000: c <= 9'b11100111;
				8'b101110: c <= 9'b110111000;
				8'b1000001: c <= 9'b110100100;
				default: c <= 9'b0;
			endcase
			9'b1011011 : case(di)
				8'b1000011: c <= 9'b111010110;
				8'b101000: c <= 9'b10111110;
				8'b111010: c <= 9'b10101110;
				8'b110110: c <= 9'b101110111;
				8'b1100100: c <= 9'b10001111;
				8'b1000000: c <= 9'b10000011;
				8'b1110110: c <= 9'b100001100;
				8'b100101: c <= 9'b100110010;
				8'b101111: c <= 9'b110111001;
				8'b100110: c <= 9'b10101001;
				8'b1100011: c <= 9'b111011001;
				8'b1001000: c <= 9'b101110111;
				8'b111000: c <= 9'b111100000;
				8'b110001: c <= 9'b101001010;
				8'b1010111: c <= 9'b111011110;
				8'b1001110: c <= 9'b101100010;
				8'b1101010: c <= 9'b100000101;
				8'b1001001: c <= 9'b10101011;
				8'b1100000: c <= 9'b11001011;
				8'b110111: c <= 9'b1100010;
				8'b1011101: c <= 9'b11011010;
				8'b1011011: c <= 9'b1000000;
				8'b111001: c <= 9'b10011011;
				8'b1001010: c <= 9'b110011010;
				8'b110011: c <= 9'b10011010;
				8'b1101100: c <= 9'b111001000;
				8'b1110111: c <= 9'b10011100;
				8'b101011: c <= 9'b110011;
				8'b1101011: c <= 9'b101001001;
				8'b111100: c <= 9'b110101010;
				8'b1000111: c <= 9'b10010;
				8'b1011111: c <= 9'b111000011;
				8'b1110100: c <= 9'b11011001;
				8'b101101: c <= 9'b10110111;
				8'b1010011: c <= 9'b110001110;
				8'b1100001: c <= 9'b100000110;
				8'b110101: c <= 9'b11000000;
				8'b1000100: c <= 9'b101010;
				8'b1010001: c <= 9'b1100100;
				8'b1010100: c <= 9'b100010;
				8'b1100110: c <= 9'b10001000;
				8'b101010: c <= 9'b111111110;
				8'b1011110: c <= 9'b110011000;
				8'b1100111: c <= 9'b101101011;
				8'b1011010: c <= 9'b10110100;
				8'b1000010: c <= 9'b1100000;
				8'b111101: c <= 9'b1000101;
				8'b110000: c <= 9'b100100101;
				8'b111110: c <= 9'b10100010;
				8'b1100010: c <= 9'b101001;
				8'b1110000: c <= 9'b10111100;
				8'b1101001: c <= 9'b100001111;
				8'b1110011: c <= 9'b1111011;
				8'b1001100: c <= 9'b101111110;
				8'b100001: c <= 9'b100011011;
				8'b1000110: c <= 9'b10;
				8'b1110010: c <= 9'b10110101;
				8'b1010000: c <= 9'b1110001;
				8'b1111010: c <= 9'b10110;
				8'b1010101: c <= 9'b110011110;
				8'b111011: c <= 9'b1001000;
				8'b1001101: c <= 9'b1011000;
				8'b111111: c <= 9'b11010;
				8'b1101110: c <= 9'b111011111;
				8'b1111011: c <= 9'b111011111;
				8'b1001011: c <= 9'b11011110;
				8'b1101111: c <= 9'b110000011;
				8'b1101000: c <= 9'b101011;
				8'b101100: c <= 9'b100110011;
				8'b100100: c <= 9'b101001000;
				8'b1111000: c <= 9'b101100100;
				8'b1000101: c <= 9'b11011110;
				8'b1011001: c <= 9'b100001110;
				8'b110100: c <= 9'b100111001;
				8'b1111001: c <= 9'b1111;
				8'b1110001: c <= 9'b111001110;
				8'b1001111: c <= 9'b10000001;
				8'b1100101: c <= 9'b10000011;
				8'b1111110: c <= 9'b11100110;
				8'b1111100: c <= 9'b11110000;
				8'b1010110: c <= 9'b1000010;
				8'b110010: c <= 9'b11110100;
				8'b1101101: c <= 9'b10001001;
				8'b100011: c <= 9'b101110100;
				8'b1110101: c <= 9'b111000000;
				8'b1111101: c <= 9'b1101100;
				8'b101001: c <= 9'b10011000;
				8'b1010010: c <= 9'b11111001;
				8'b1011000: c <= 9'b110010011;
				8'b101110: c <= 9'b10111100;
				8'b1000001: c <= 9'b11100110;
				default: c <= 9'b0;
			endcase
			9'b100101110 : case(di)
				8'b1000011: c <= 9'b110000010;
				8'b101000: c <= 9'b101100100;
				8'b111010: c <= 9'b1100011;
				8'b110110: c <= 9'b10110010;
				8'b1100100: c <= 9'b101111110;
				8'b1000000: c <= 9'b110001011;
				8'b1110110: c <= 9'b110110100;
				8'b100101: c <= 9'b100001111;
				8'b101111: c <= 9'b1000111;
				8'b100110: c <= 9'b11110100;
				8'b1100011: c <= 9'b101101001;
				8'b1001000: c <= 9'b100010;
				8'b111000: c <= 9'b100101000;
				8'b110001: c <= 9'b111000;
				8'b1010111: c <= 9'b10000;
				8'b1001110: c <= 9'b100010;
				8'b1101010: c <= 9'b11011000;
				8'b1001001: c <= 9'b110100110;
				8'b1100000: c <= 9'b101111000;
				8'b110111: c <= 9'b10010000;
				8'b1011101: c <= 9'b101011101;
				8'b1011011: c <= 9'b110100111;
				8'b111001: c <= 9'b100010000;
				8'b1001010: c <= 9'b101010100;
				8'b110011: c <= 9'b111111111;
				8'b1101100: c <= 9'b110001;
				8'b1110111: c <= 9'b101100000;
				8'b101011: c <= 9'b110000;
				8'b1101011: c <= 9'b100101;
				8'b111100: c <= 9'b10110101;
				8'b1000111: c <= 9'b1011;
				8'b1011111: c <= 9'b111000110;
				8'b1110100: c <= 9'b111001111;
				8'b101101: c <= 9'b11010111;
				8'b1010011: c <= 9'b10010111;
				8'b1100001: c <= 9'b10101000;
				8'b110101: c <= 9'b100011011;
				8'b1000100: c <= 9'b11010001;
				8'b1010001: c <= 9'b10001110;
				8'b1010100: c <= 9'b11001000;
				8'b1100110: c <= 9'b100110;
				8'b101010: c <= 9'b100101010;
				8'b1011110: c <= 9'b10101;
				8'b1100111: c <= 9'b111110011;
				8'b1011010: c <= 9'b111000100;
				8'b1000010: c <= 9'b100000000;
				8'b111101: c <= 9'b111000000;
				8'b110000: c <= 9'b111100;
				8'b111110: c <= 9'b11001001;
				8'b1100010: c <= 9'b11011000;
				8'b1110000: c <= 9'b11111001;
				8'b1101001: c <= 9'b11111110;
				8'b1110011: c <= 9'b1001010;
				8'b1001100: c <= 9'b111000010;
				8'b100001: c <= 9'b10001000;
				8'b1000110: c <= 9'b1010101;
				8'b1110010: c <= 9'b111101001;
				8'b1010000: c <= 9'b11100000;
				8'b1111010: c <= 9'b1001111;
				8'b1010101: c <= 9'b111011011;
				8'b111011: c <= 9'b10010100;
				8'b1001101: c <= 9'b110011000;
				8'b111111: c <= 9'b10110110;
				8'b1101110: c <= 9'b110011101;
				8'b1111011: c <= 9'b1110001;
				8'b1001011: c <= 9'b111001111;
				8'b1101111: c <= 9'b111100010;
				8'b1101000: c <= 9'b101110011;
				8'b101100: c <= 9'b101111001;
				8'b100100: c <= 9'b10111000;
				8'b1111000: c <= 9'b100101010;
				8'b1000101: c <= 9'b10100101;
				8'b1011001: c <= 9'b110010111;
				8'b110100: c <= 9'b110100111;
				8'b1111001: c <= 9'b101001001;
				8'b1110001: c <= 9'b100001001;
				8'b1001111: c <= 9'b110110100;
				8'b1100101: c <= 9'b110100101;
				8'b1111110: c <= 9'b100101011;
				8'b1111100: c <= 9'b101010010;
				8'b1010110: c <= 9'b100010011;
				8'b110010: c <= 9'b110001010;
				8'b1101101: c <= 9'b101110010;
				8'b100011: c <= 9'b111000010;
				8'b1110101: c <= 9'b100001;
				8'b1111101: c <= 9'b111001001;
				8'b101001: c <= 9'b110101110;
				8'b1010010: c <= 9'b111011010;
				8'b1011000: c <= 9'b111000110;
				8'b101110: c <= 9'b1011000;
				8'b1000001: c <= 9'b100000100;
				default: c <= 9'b0;
			endcase
			9'b110011110 : case(di)
				8'b1000011: c <= 9'b101001001;
				8'b101000: c <= 9'b10001111;
				8'b111010: c <= 9'b110011;
				8'b110110: c <= 9'b101001001;
				8'b1100100: c <= 9'b111000000;
				8'b1000000: c <= 9'b1011011;
				8'b1110110: c <= 9'b11100111;
				8'b100101: c <= 9'b110100000;
				8'b101111: c <= 9'b11000001;
				8'b100110: c <= 9'b111110110;
				8'b1100011: c <= 9'b11111110;
				8'b1001000: c <= 9'b110010010;
				8'b111000: c <= 9'b100110000;
				8'b110001: c <= 9'b100000101;
				8'b1010111: c <= 9'b111011111;
				8'b1001110: c <= 9'b100111011;
				8'b1101010: c <= 9'b111101010;
				8'b1001001: c <= 9'b11010011;
				8'b1100000: c <= 9'b100111;
				8'b110111: c <= 9'b10001111;
				8'b1011101: c <= 9'b11010101;
				8'b1011011: c <= 9'b110101010;
				8'b111001: c <= 9'b111010;
				8'b1001010: c <= 9'b11100;
				8'b110011: c <= 9'b100011100;
				8'b1101100: c <= 9'b1110;
				8'b1110111: c <= 9'b11101100;
				8'b101011: c <= 9'b111100;
				8'b1101011: c <= 9'b101010111;
				8'b111100: c <= 9'b1010010;
				8'b1000111: c <= 9'b11100;
				8'b1011111: c <= 9'b1001000;
				8'b1110100: c <= 9'b111100000;
				8'b101101: c <= 9'b110001000;
				8'b1010011: c <= 9'b101011000;
				8'b1100001: c <= 9'b1000011;
				8'b110101: c <= 9'b1111110;
				8'b1000100: c <= 9'b10111100;
				8'b1010001: c <= 9'b100110110;
				8'b1010100: c <= 9'b111;
				8'b1100110: c <= 9'b111100101;
				8'b101010: c <= 9'b11101101;
				8'b1011110: c <= 9'b100100110;
				8'b1100111: c <= 9'b1101110;
				8'b1011010: c <= 9'b11;
				8'b1000010: c <= 9'b110110100;
				8'b111101: c <= 9'b101101011;
				8'b110000: c <= 9'b111101001;
				8'b111110: c <= 9'b11001101;
				8'b1100010: c <= 9'b100101;
				8'b1110000: c <= 9'b111100001;
				8'b1101001: c <= 9'b110011110;
				8'b1110011: c <= 9'b101111010;
				8'b1001100: c <= 9'b11011100;
				8'b100001: c <= 9'b110000111;
				8'b1000110: c <= 9'b10010100;
				8'b1110010: c <= 9'b1110100;
				8'b1010000: c <= 9'b1100;
				8'b1111010: c <= 9'b1010101;
				8'b1010101: c <= 9'b11100101;
				8'b111011: c <= 9'b11110;
				8'b1001101: c <= 9'b111101010;
				8'b111111: c <= 9'b110011;
				8'b1101110: c <= 9'b11001;
				8'b1111011: c <= 9'b11000;
				8'b1001011: c <= 9'b110011010;
				8'b1101111: c <= 9'b1010111;
				8'b1101000: c <= 9'b11111100;
				8'b101100: c <= 9'b10011001;
				8'b100100: c <= 9'b100110110;
				8'b1111000: c <= 9'b1001000;
				8'b1000101: c <= 9'b100011111;
				8'b1011001: c <= 9'b111010111;
				8'b110100: c <= 9'b100100111;
				8'b1111001: c <= 9'b1111010;
				8'b1110001: c <= 9'b1110010;
				8'b1001111: c <= 9'b1100000;
				8'b1100101: c <= 9'b100101100;
				8'b1111110: c <= 9'b110100101;
				8'b1111100: c <= 9'b10010001;
				8'b1010110: c <= 9'b110111110;
				8'b110010: c <= 9'b11010000;
				8'b1101101: c <= 9'b11001100;
				8'b100011: c <= 9'b110010;
				8'b1110101: c <= 9'b111111;
				8'b1111101: c <= 9'b11010000;
				8'b101001: c <= 9'b101100110;
				8'b1010010: c <= 9'b1110011;
				8'b1011000: c <= 9'b100001;
				8'b101110: c <= 9'b111100101;
				8'b1000001: c <= 9'b10110110;
				default: c <= 9'b0;
			endcase
			9'b110001010 : case(di)
				8'b1000011: c <= 9'b101010111;
				8'b101000: c <= 9'b101001000;
				8'b111010: c <= 9'b10010011;
				8'b110110: c <= 9'b101010001;
				8'b1100100: c <= 9'b101001010;
				8'b1000000: c <= 9'b110110100;
				8'b1110110: c <= 9'b111101;
				8'b100101: c <= 9'b10;
				8'b101111: c <= 9'b10010;
				8'b100110: c <= 9'b111011101;
				8'b1100011: c <= 9'b10010000;
				8'b1001000: c <= 9'b11000001;
				8'b111000: c <= 9'b10111111;
				8'b110001: c <= 9'b100100001;
				8'b1010111: c <= 9'b110001110;
				8'b1001110: c <= 9'b1000111;
				8'b1101010: c <= 9'b100010011;
				8'b1001001: c <= 9'b110000111;
				8'b1100000: c <= 9'b110110011;
				8'b110111: c <= 9'b110111011;
				8'b1011101: c <= 9'b1011001;
				8'b1011011: c <= 9'b10100011;
				8'b111001: c <= 9'b11110001;
				8'b1001010: c <= 9'b1001111;
				8'b110011: c <= 9'b110011110;
				8'b1101100: c <= 9'b11010001;
				8'b1110111: c <= 9'b111010100;
				8'b101011: c <= 9'b101111111;
				8'b1101011: c <= 9'b1100100;
				8'b111100: c <= 9'b110000010;
				8'b1000111: c <= 9'b100001100;
				8'b1011111: c <= 9'b1100;
				8'b1110100: c <= 9'b100111110;
				8'b101101: c <= 9'b101100101;
				8'b1010011: c <= 9'b111100110;
				8'b1100001: c <= 9'b101110110;
				8'b110101: c <= 9'b1100011;
				8'b1000100: c <= 9'b10110;
				8'b1010001: c <= 9'b111110110;
				8'b1010100: c <= 9'b110000111;
				8'b1100110: c <= 9'b10110001;
				8'b101010: c <= 9'b10101;
				8'b1011110: c <= 9'b1101001;
				8'b1100111: c <= 9'b111111001;
				8'b1011010: c <= 9'b110111100;
				8'b1000010: c <= 9'b10100100;
				8'b111101: c <= 9'b1;
				8'b110000: c <= 9'b1001100;
				8'b111110: c <= 9'b101111111;
				8'b1100010: c <= 9'b101010101;
				8'b1110000: c <= 9'b100100001;
				8'b1101001: c <= 9'b100111110;
				8'b1110011: c <= 9'b1110100;
				8'b1001100: c <= 9'b11000110;
				8'b100001: c <= 9'b1100110;
				8'b1000110: c <= 9'b100000110;
				8'b1110010: c <= 9'b110001011;
				8'b1010000: c <= 9'b100010001;
				8'b1111010: c <= 9'b101101001;
				8'b1010101: c <= 9'b100010101;
				8'b111011: c <= 9'b101110010;
				8'b1001101: c <= 9'b10110;
				8'b111111: c <= 9'b11010;
				8'b1101110: c <= 9'b1111001;
				8'b1111011: c <= 9'b100101110;
				8'b1001011: c <= 9'b110110011;
				8'b1101111: c <= 9'b111001011;
				8'b1101000: c <= 9'b111001111;
				8'b101100: c <= 9'b110110100;
				8'b100100: c <= 9'b1010101;
				8'b1111000: c <= 9'b11110100;
				8'b1000101: c <= 9'b110100110;
				8'b1011001: c <= 9'b101010111;
				8'b110100: c <= 9'b10101;
				8'b1111001: c <= 9'b1001001;
				8'b1110001: c <= 9'b1001001;
				8'b1001111: c <= 9'b100001100;
				8'b1100101: c <= 9'b1001100;
				8'b1111110: c <= 9'b101110011;
				8'b1111100: c <= 9'b11011110;
				8'b1010110: c <= 9'b111010010;
				8'b110010: c <= 9'b10111101;
				8'b1101101: c <= 9'b110000001;
				8'b100011: c <= 9'b110110010;
				8'b1110101: c <= 9'b110110010;
				8'b1111101: c <= 9'b100010001;
				8'b101001: c <= 9'b10011101;
				8'b1010010: c <= 9'b1001010;
				8'b1011000: c <= 9'b1110111;
				8'b101110: c <= 9'b1101000;
				8'b1000001: c <= 9'b110000110;
				default: c <= 9'b0;
			endcase
			9'b110011011 : case(di)
				8'b1000011: c <= 9'b10101101;
				8'b101000: c <= 9'b11110001;
				8'b111010: c <= 9'b11000000;
				8'b110110: c <= 9'b101011011;
				8'b1100100: c <= 9'b11001111;
				8'b1000000: c <= 9'b1111100;
				8'b1110110: c <= 9'b10110;
				8'b100101: c <= 9'b11000010;
				8'b101111: c <= 9'b111001011;
				8'b100110: c <= 9'b101000100;
				8'b1100011: c <= 9'b111111001;
				8'b1001000: c <= 9'b100000111;
				8'b111000: c <= 9'b1010101;
				8'b110001: c <= 9'b100100110;
				8'b1010111: c <= 9'b10000101;
				8'b1001110: c <= 9'b11111100;
				8'b1101010: c <= 9'b11001000;
				8'b1001001: c <= 9'b101010101;
				8'b1100000: c <= 9'b101;
				8'b110111: c <= 9'b10000010;
				8'b1011101: c <= 9'b100001010;
				8'b1011011: c <= 9'b111001110;
				8'b111001: c <= 9'b1101;
				8'b1001010: c <= 9'b100110;
				8'b110011: c <= 9'b100101010;
				8'b1101100: c <= 9'b101100110;
				8'b1110111: c <= 9'b1100101;
				8'b101011: c <= 9'b100100000;
				8'b1101011: c <= 9'b110000011;
				8'b111100: c <= 9'b11111101;
				8'b1000111: c <= 9'b101011110;
				8'b1011111: c <= 9'b110110;
				8'b1110100: c <= 9'b100001110;
				8'b101101: c <= 9'b111101001;
				8'b1010011: c <= 9'b101111111;
				8'b1100001: c <= 9'b100;
				8'b110101: c <= 9'b11100110;
				8'b1000100: c <= 9'b111101001;
				8'b1010001: c <= 9'b10111000;
				8'b1010100: c <= 9'b111100110;
				8'b1100110: c <= 9'b101011111;
				8'b101010: c <= 9'b10001011;
				8'b1011110: c <= 9'b11101111;
				8'b1100111: c <= 9'b110010010;
				8'b1011010: c <= 9'b111001;
				8'b1000010: c <= 9'b1001111;
				8'b111101: c <= 9'b110101111;
				8'b110000: c <= 9'b100001;
				8'b111110: c <= 9'b1010000;
				8'b1100010: c <= 9'b11111110;
				8'b1110000: c <= 9'b111101101;
				8'b1101001: c <= 9'b110001000;
				8'b1110011: c <= 9'b111111111;
				8'b1001100: c <= 9'b10001110;
				8'b100001: c <= 9'b10111001;
				8'b1000110: c <= 9'b110111110;
				8'b1110010: c <= 9'b10000011;
				8'b1010000: c <= 9'b11010001;
				8'b1111010: c <= 9'b11001110;
				8'b1010101: c <= 9'b110110010;
				8'b111011: c <= 9'b111111101;
				8'b1001101: c <= 9'b101000001;
				8'b111111: c <= 9'b110111100;
				8'b1101110: c <= 9'b101100001;
				8'b1111011: c <= 9'b110011110;
				8'b1001011: c <= 9'b11100000;
				8'b1101111: c <= 9'b111011011;
				8'b1101000: c <= 9'b110100011;
				8'b101100: c <= 9'b1010111;
				8'b100100: c <= 9'b111001001;
				8'b1111000: c <= 9'b110110011;
				8'b1000101: c <= 9'b1000010;
				8'b1011001: c <= 9'b11110010;
				8'b110100: c <= 9'b11000010;
				8'b1111001: c <= 9'b100011001;
				8'b1110001: c <= 9'b10101110;
				8'b1001111: c <= 9'b1100010;
				8'b1100101: c <= 9'b11110001;
				8'b1111110: c <= 9'b11110101;
				8'b1111100: c <= 9'b110011;
				8'b1010110: c <= 9'b11001111;
				8'b110010: c <= 9'b110001011;
				8'b1101101: c <= 9'b11000111;
				8'b100011: c <= 9'b111110000;
				8'b1110101: c <= 9'b101110110;
				8'b1111101: c <= 9'b10001100;
				8'b101001: c <= 9'b100101010;
				8'b1010010: c <= 9'b100010;
				8'b1011000: c <= 9'b1000110;
				8'b101110: c <= 9'b1110001;
				8'b1000001: c <= 9'b101101110;
				default: c <= 9'b0;
			endcase
			9'b1111010 : case(di)
				8'b1000011: c <= 9'b100111110;
				8'b101000: c <= 9'b100011111;
				8'b111010: c <= 9'b101110101;
				8'b110110: c <= 9'b1101010;
				8'b1100100: c <= 9'b100100000;
				8'b1000000: c <= 9'b1001;
				8'b1110110: c <= 9'b100011111;
				8'b100101: c <= 9'b10101;
				8'b101111: c <= 9'b1010110;
				8'b100110: c <= 9'b10100011;
				8'b1100011: c <= 9'b1110101;
				8'b1001000: c <= 9'b10101110;
				8'b111000: c <= 9'b111100000;
				8'b110001: c <= 9'b101000111;
				8'b1010111: c <= 9'b101101110;
				8'b1001110: c <= 9'b1000101;
				8'b1101010: c <= 9'b101010011;
				8'b1001001: c <= 9'b100111;
				8'b1100000: c <= 9'b1111010;
				8'b110111: c <= 9'b111111111;
				8'b1011101: c <= 9'b111000101;
				8'b1011011: c <= 9'b101010010;
				8'b111001: c <= 9'b100100011;
				8'b1001010: c <= 9'b11010000;
				8'b110011: c <= 9'b111010000;
				8'b1101100: c <= 9'b100101010;
				8'b1110111: c <= 9'b10110011;
				8'b101011: c <= 9'b1100;
				8'b1101011: c <= 9'b11000110;
				8'b111100: c <= 9'b11000100;
				8'b1000111: c <= 9'b1000111;
				8'b1011111: c <= 9'b110001110;
				8'b1110100: c <= 9'b11010010;
				8'b101101: c <= 9'b101100111;
				8'b1010011: c <= 9'b100000000;
				8'b1100001: c <= 9'b10110010;
				8'b110101: c <= 9'b101010111;
				8'b1000100: c <= 9'b11111001;
				8'b1010001: c <= 9'b1010110;
				8'b1010100: c <= 9'b100000000;
				8'b1100110: c <= 9'b110100111;
				8'b101010: c <= 9'b100111010;
				8'b1011110: c <= 9'b11100000;
				8'b1100111: c <= 9'b100101110;
				8'b1011010: c <= 9'b101101011;
				8'b1000010: c <= 9'b111100111;
				8'b111101: c <= 9'b111011100;
				8'b110000: c <= 9'b11111000;
				8'b111110: c <= 9'b1101101;
				8'b1100010: c <= 9'b100101001;
				8'b1110000: c <= 9'b1011100;
				8'b1101001: c <= 9'b111011111;
				8'b1110011: c <= 9'b1001011;
				8'b1001100: c <= 9'b101111000;
				8'b100001: c <= 9'b1101100;
				8'b1000110: c <= 9'b11001010;
				8'b1110010: c <= 9'b11001010;
				8'b1010000: c <= 9'b11011;
				8'b1111010: c <= 9'b1010000;
				8'b1010101: c <= 9'b10011101;
				8'b111011: c <= 9'b110010100;
				8'b1001101: c <= 9'b1100011;
				8'b111111: c <= 9'b10011;
				8'b1101110: c <= 9'b100010111;
				8'b1111011: c <= 9'b10111100;
				8'b1001011: c <= 9'b10101011;
				8'b1101111: c <= 9'b110001100;
				8'b1101000: c <= 9'b101110011;
				8'b101100: c <= 9'b1000001;
				8'b100100: c <= 9'b110011;
				8'b1111000: c <= 9'b100000100;
				8'b1000101: c <= 9'b1000010;
				8'b1011001: c <= 9'b111000;
				8'b110100: c <= 9'b11100010;
				8'b1111001: c <= 9'b110111110;
				8'b1110001: c <= 9'b110101001;
				8'b1001111: c <= 9'b101001010;
				8'b1100101: c <= 9'b110100011;
				8'b1111110: c <= 9'b101100111;
				8'b1111100: c <= 9'b10101110;
				8'b1010110: c <= 9'b1001100;
				8'b110010: c <= 9'b1100;
				8'b1101101: c <= 9'b10100100;
				8'b100011: c <= 9'b10101110;
				8'b1110101: c <= 9'b11111010;
				8'b1111101: c <= 9'b110011100;
				8'b101001: c <= 9'b101110110;
				8'b1010010: c <= 9'b1101101;
				8'b1011000: c <= 9'b110101011;
				8'b101110: c <= 9'b1101001;
				8'b1000001: c <= 9'b100011001;
				default: c <= 9'b0;
			endcase
			9'b1001110 : case(di)
				8'b1000011: c <= 9'b101011001;
				8'b101000: c <= 9'b1110100;
				8'b111010: c <= 9'b110010010;
				8'b110110: c <= 9'b100110;
				8'b1100100: c <= 9'b10110100;
				8'b1000000: c <= 9'b111000;
				8'b1110110: c <= 9'b11001100;
				8'b100101: c <= 9'b101101011;
				8'b101111: c <= 9'b11;
				8'b100110: c <= 9'b101101101;
				8'b1100011: c <= 9'b1100000;
				8'b1001000: c <= 9'b111111;
				8'b111000: c <= 9'b101000110;
				8'b110001: c <= 9'b101011111;
				8'b1010111: c <= 9'b1111001;
				8'b1001110: c <= 9'b101110111;
				8'b1101010: c <= 9'b101110101;
				8'b1001001: c <= 9'b11100101;
				8'b1100000: c <= 9'b100111;
				8'b110111: c <= 9'b100000001;
				8'b1011101: c <= 9'b11110001;
				8'b1011011: c <= 9'b101111001;
				8'b111001: c <= 9'b1110101;
				8'b1001010: c <= 9'b100111110;
				8'b110011: c <= 9'b100110000;
				8'b1101100: c <= 9'b10001001;
				8'b1110111: c <= 9'b100011011;
				8'b101011: c <= 9'b100001111;
				8'b1101011: c <= 9'b10000000;
				8'b111100: c <= 9'b101111000;
				8'b1000111: c <= 9'b111000111;
				8'b1011111: c <= 9'b101101011;
				8'b1110100: c <= 9'b1111;
				8'b101101: c <= 9'b100111010;
				8'b1010011: c <= 9'b10;
				8'b1100001: c <= 9'b1001111;
				8'b110101: c <= 9'b1001111;
				8'b1000100: c <= 9'b11011100;
				8'b1010001: c <= 9'b11001111;
				8'b1010100: c <= 9'b100100001;
				8'b1100110: c <= 9'b1010110;
				8'b101010: c <= 9'b1101110;
				8'b1011110: c <= 9'b110011;
				8'b1100111: c <= 9'b10101010;
				8'b1011010: c <= 9'b110010010;
				8'b1000010: c <= 9'b10100;
				8'b111101: c <= 9'b100011010;
				8'b110000: c <= 9'b11110000;
				8'b111110: c <= 9'b11110000;
				8'b1100010: c <= 9'b1100110;
				8'b1110000: c <= 9'b111100110;
				8'b1101001: c <= 9'b111011010;
				8'b1110011: c <= 9'b11010101;
				8'b1001100: c <= 9'b1000011;
				8'b100001: c <= 9'b11110111;
				8'b1000110: c <= 9'b101110;
				8'b1110010: c <= 9'b111100001;
				8'b1010000: c <= 9'b1010001;
				8'b1111010: c <= 9'b100011000;
				8'b1010101: c <= 9'b100011111;
				8'b111011: c <= 9'b100010010;
				8'b1001101: c <= 9'b11111100;
				8'b111111: c <= 9'b1010011;
				8'b1101110: c <= 9'b11010010;
				8'b1111011: c <= 9'b101000111;
				8'b1001011: c <= 9'b10101100;
				8'b1101111: c <= 9'b1010101;
				8'b1101000: c <= 9'b110010010;
				8'b101100: c <= 9'b100111101;
				8'b100100: c <= 9'b111100100;
				8'b1111000: c <= 9'b1000101;
				8'b1000101: c <= 9'b10101000;
				8'b1011001: c <= 9'b10001101;
				8'b110100: c <= 9'b1101110;
				8'b1111001: c <= 9'b101000001;
				8'b1110001: c <= 9'b10110110;
				8'b1001111: c <= 9'b101010101;
				8'b1100101: c <= 9'b100100001;
				8'b1111110: c <= 9'b110000011;
				8'b1111100: c <= 9'b11010111;
				8'b1010110: c <= 9'b110000101;
				8'b110010: c <= 9'b10111101;
				8'b1101101: c <= 9'b11001010;
				8'b100011: c <= 9'b100101110;
				8'b1110101: c <= 9'b110001000;
				8'b1111101: c <= 9'b110111;
				8'b101001: c <= 9'b10110011;
				8'b1010010: c <= 9'b111111110;
				8'b1011000: c <= 9'b111101110;
				8'b101110: c <= 9'b11001110;
				8'b1000001: c <= 9'b1101101;
				default: c <= 9'b0;
			endcase
			9'b101011011 : case(di)
				8'b1000011: c <= 9'b10000011;
				8'b101000: c <= 9'b11100110;
				8'b111010: c <= 9'b110001101;
				8'b110110: c <= 9'b111011001;
				8'b1100100: c <= 9'b11010011;
				8'b1000000: c <= 9'b11011000;
				8'b1110110: c <= 9'b111010001;
				8'b100101: c <= 9'b11001100;
				8'b101111: c <= 9'b10001101;
				8'b100110: c <= 9'b1111100;
				8'b1100011: c <= 9'b110111100;
				8'b1001000: c <= 9'b100101100;
				8'b111000: c <= 9'b11100110;
				8'b110001: c <= 9'b11000000;
				8'b1010111: c <= 9'b10100010;
				8'b1001110: c <= 9'b10111110;
				8'b1101010: c <= 9'b110001111;
				8'b1001001: c <= 9'b1010001;
				8'b1100000: c <= 9'b11;
				8'b110111: c <= 9'b110011111;
				8'b1011101: c <= 9'b111011111;
				8'b1011011: c <= 9'b101000011;
				8'b111001: c <= 9'b100010;
				8'b1001010: c <= 9'b1111110;
				8'b110011: c <= 9'b1001;
				8'b1101100: c <= 9'b11100100;
				8'b1110111: c <= 9'b1111110;
				8'b101011: c <= 9'b1001001;
				8'b1101011: c <= 9'b11101111;
				8'b111100: c <= 9'b100110111;
				8'b1000111: c <= 9'b111111000;
				8'b1011111: c <= 9'b1100111;
				8'b1110100: c <= 9'b1101110;
				8'b101101: c <= 9'b11000000;
				8'b1010011: c <= 9'b110111100;
				8'b1100001: c <= 9'b11010101;
				8'b110101: c <= 9'b11011110;
				8'b1000100: c <= 9'b110111011;
				8'b1010001: c <= 9'b10111001;
				8'b1010100: c <= 9'b10011000;
				8'b1100110: c <= 9'b10000110;
				8'b101010: c <= 9'b10101101;
				8'b1011110: c <= 9'b110100011;
				8'b1100111: c <= 9'b10101010;
				8'b1011010: c <= 9'b1100100;
				8'b1000010: c <= 9'b111;
				8'b111101: c <= 9'b110010101;
				8'b110000: c <= 9'b11101100;
				8'b111110: c <= 9'b10110110;
				8'b1100010: c <= 9'b11011000;
				8'b1110000: c <= 9'b10000111;
				8'b1101001: c <= 9'b111001001;
				8'b1110011: c <= 9'b100111000;
				8'b1001100: c <= 9'b110000111;
				8'b100001: c <= 9'b100101000;
				8'b1000110: c <= 9'b101011010;
				8'b1110010: c <= 9'b110100110;
				8'b1010000: c <= 9'b1001110;
				8'b1111010: c <= 9'b11001010;
				8'b1010101: c <= 9'b101101111;
				8'b111011: c <= 9'b10110011;
				8'b1001101: c <= 9'b1000000;
				8'b111111: c <= 9'b11110;
				8'b1101110: c <= 9'b10011000;
				8'b1111011: c <= 9'b101101111;
				8'b1001011: c <= 9'b10100011;
				8'b1101111: c <= 9'b110001001;
				8'b1101000: c <= 9'b1010000;
				8'b101100: c <= 9'b11110110;
				8'b100100: c <= 9'b11100100;
				8'b1111000: c <= 9'b1001100;
				8'b1000101: c <= 9'b1110011;
				8'b1011001: c <= 9'b1001101;
				8'b110100: c <= 9'b110010101;
				8'b1111001: c <= 9'b10111100;
				8'b1110001: c <= 9'b1111011;
				8'b1001111: c <= 9'b1101110;
				8'b1100101: c <= 9'b110100001;
				8'b1111110: c <= 9'b11011000;
				8'b1111100: c <= 9'b110101111;
				8'b1010110: c <= 9'b111101101;
				8'b110010: c <= 9'b111001000;
				8'b1101101: c <= 9'b1011111;
				8'b100011: c <= 9'b10010;
				8'b1110101: c <= 9'b11011110;
				8'b1111101: c <= 9'b110110;
				8'b101001: c <= 9'b110111100;
				8'b1010010: c <= 9'b10110100;
				8'b1011000: c <= 9'b110010011;
				8'b101110: c <= 9'b10001010;
				8'b1000001: c <= 9'b110111010;
				default: c <= 9'b0;
			endcase
			9'b10011101 : case(di)
				8'b1000011: c <= 9'b110100111;
				8'b101000: c <= 9'b10111110;
				8'b111010: c <= 9'b10001101;
				8'b110110: c <= 9'b100101;
				8'b1100100: c <= 9'b101100100;
				8'b1000000: c <= 9'b11001010;
				8'b1110110: c <= 9'b10000010;
				8'b100101: c <= 9'b1;
				8'b101111: c <= 9'b101010110;
				8'b100110: c <= 9'b101100;
				8'b1100011: c <= 9'b101101010;
				8'b1001000: c <= 9'b10010111;
				8'b111000: c <= 9'b101101011;
				8'b110001: c <= 9'b111111010;
				8'b1010111: c <= 9'b1100111;
				8'b1001110: c <= 9'b100100;
				8'b1101010: c <= 9'b110110111;
				8'b1001001: c <= 9'b111110110;
				8'b1100000: c <= 9'b111100001;
				8'b110111: c <= 9'b111010110;
				8'b1011101: c <= 9'b100000011;
				8'b1011011: c <= 9'b11110000;
				8'b111001: c <= 9'b1100111;
				8'b1001010: c <= 9'b110010111;
				8'b110011: c <= 9'b1011011;
				8'b1101100: c <= 9'b111001110;
				8'b1110111: c <= 9'b10010100;
				8'b101011: c <= 9'b11001111;
				8'b1101011: c <= 9'b111;
				8'b111100: c <= 9'b111111110;
				8'b1000111: c <= 9'b111000111;
				8'b1011111: c <= 9'b110001110;
				8'b1110100: c <= 9'b101;
				8'b101101: c <= 9'b101101110;
				8'b1010011: c <= 9'b1000110;
				8'b1100001: c <= 9'b1000011;
				8'b110101: c <= 9'b100011111;
				8'b1000100: c <= 9'b10110111;
				8'b1010001: c <= 9'b100111001;
				8'b1010100: c <= 9'b101001000;
				8'b1100110: c <= 9'b11111110;
				8'b101010: c <= 9'b1111011;
				8'b1011110: c <= 9'b101001110;
				8'b1100111: c <= 9'b1011;
				8'b1011010: c <= 9'b101010110;
				8'b1000010: c <= 9'b110011110;
				8'b111101: c <= 9'b110010001;
				8'b110000: c <= 9'b10;
				8'b111110: c <= 9'b11101011;
				8'b1100010: c <= 9'b11011010;
				8'b1110000: c <= 9'b10110110;
				8'b1101001: c <= 9'b10100;
				8'b1110011: c <= 9'b11011110;
				8'b1001100: c <= 9'b101010111;
				8'b100001: c <= 9'b100001011;
				8'b1000110: c <= 9'b111000000;
				8'b1110010: c <= 9'b111001110;
				8'b1010000: c <= 9'b101011010;
				8'b1111010: c <= 9'b10011001;
				8'b1010101: c <= 9'b111000000;
				8'b111011: c <= 9'b100011011;
				8'b1001101: c <= 9'b111011100;
				8'b111111: c <= 9'b10110110;
				8'b1101110: c <= 9'b10101011;
				8'b1111011: c <= 9'b11000000;
				8'b1001011: c <= 9'b111101111;
				8'b1101111: c <= 9'b101011010;
				8'b1101000: c <= 9'b110011101;
				8'b101100: c <= 9'b11111001;
				8'b100100: c <= 9'b101000110;
				8'b1111000: c <= 9'b1001;
				8'b1000101: c <= 9'b11111;
				8'b1011001: c <= 9'b11001100;
				8'b110100: c <= 9'b101000111;
				8'b1111001: c <= 9'b101100110;
				8'b1110001: c <= 9'b111000010;
				8'b1001111: c <= 9'b11000111;
				8'b1100101: c <= 9'b100011000;
				8'b1111110: c <= 9'b100100001;
				8'b1111100: c <= 9'b110111010;
				8'b1010110: c <= 9'b111001001;
				8'b110010: c <= 9'b1011111;
				8'b1101101: c <= 9'b10101;
				8'b100011: c <= 9'b111101001;
				8'b1110101: c <= 9'b1010101;
				8'b1111101: c <= 9'b110111100;
				8'b101001: c <= 9'b110111000;
				8'b1010010: c <= 9'b11100111;
				8'b1011000: c <= 9'b111101000;
				8'b101110: c <= 9'b111111011;
				8'b1000001: c <= 9'b10001100;
				default: c <= 9'b0;
			endcase
			9'b1010110 : case(di)
				8'b1000011: c <= 9'b10011101;
				8'b101000: c <= 9'b1011010;
				8'b111010: c <= 9'b111011101;
				8'b110110: c <= 9'b100101000;
				8'b1100100: c <= 9'b100111;
				8'b1000000: c <= 9'b11111;
				8'b1110110: c <= 9'b1011001;
				8'b100101: c <= 9'b10000011;
				8'b101111: c <= 9'b10100010;
				8'b100110: c <= 9'b1001010;
				8'b1100011: c <= 9'b110001001;
				8'b1001000: c <= 9'b10100111;
				8'b111000: c <= 9'b111110011;
				8'b110001: c <= 9'b10000011;
				8'b1010111: c <= 9'b11001100;
				8'b1001110: c <= 9'b101011110;
				8'b1101010: c <= 9'b100011100;
				8'b1001001: c <= 9'b10111011;
				8'b1100000: c <= 9'b11011001;
				8'b110111: c <= 9'b100111000;
				8'b1011101: c <= 9'b100111001;
				8'b1011011: c <= 9'b11101111;
				8'b111001: c <= 9'b11010;
				8'b1001010: c <= 9'b11110101;
				8'b110011: c <= 9'b11111011;
				8'b1101100: c <= 9'b10;
				8'b1110111: c <= 9'b1100010;
				8'b101011: c <= 9'b100011011;
				8'b1101011: c <= 9'b110000110;
				8'b111100: c <= 9'b100101;
				8'b1000111: c <= 9'b101100111;
				8'b1011111: c <= 9'b101000001;
				8'b1110100: c <= 9'b111000010;
				8'b101101: c <= 9'b101100101;
				8'b1010011: c <= 9'b10100110;
				8'b1100001: c <= 9'b11001101;
				8'b110101: c <= 9'b11000011;
				8'b1000100: c <= 9'b110100111;
				8'b1010001: c <= 9'b110111000;
				8'b1010100: c <= 9'b1111;
				8'b1100110: c <= 9'b11111011;
				8'b101010: c <= 9'b10101110;
				8'b1011110: c <= 9'b10111110;
				8'b1100111: c <= 9'b1100000;
				8'b1011010: c <= 9'b1001000;
				8'b1000010: c <= 9'b110111011;
				8'b111101: c <= 9'b1101111;
				8'b110000: c <= 9'b110101110;
				8'b111110: c <= 9'b101010100;
				8'b1100010: c <= 9'b110101110;
				8'b1110000: c <= 9'b11010101;
				8'b1101001: c <= 9'b10110111;
				8'b1110011: c <= 9'b111011100;
				8'b1001100: c <= 9'b100011111;
				8'b100001: c <= 9'b10110010;
				8'b1000110: c <= 9'b110101110;
				8'b1110010: c <= 9'b10011100;
				8'b1010000: c <= 9'b111111001;
				8'b1111010: c <= 9'b100110011;
				8'b1010101: c <= 9'b10001101;
				8'b111011: c <= 9'b100100000;
				8'b1001101: c <= 9'b110010100;
				8'b111111: c <= 9'b100101010;
				8'b1101110: c <= 9'b111111010;
				8'b1111011: c <= 9'b111100110;
				8'b1001011: c <= 9'b111001;
				8'b1101111: c <= 9'b111100;
				8'b1101000: c <= 9'b110011000;
				8'b101100: c <= 9'b100001011;
				8'b100100: c <= 9'b100000001;
				8'b1111000: c <= 9'b10111111;
				8'b1000101: c <= 9'b1011;
				8'b1011001: c <= 9'b100000000;
				8'b110100: c <= 9'b10100;
				8'b1111001: c <= 9'b101011111;
				8'b1110001: c <= 9'b10110100;
				8'b1001111: c <= 9'b100000011;
				8'b1100101: c <= 9'b101000010;
				8'b1111110: c <= 9'b110100011;
				8'b1111100: c <= 9'b11101001;
				8'b1010110: c <= 9'b110011001;
				8'b110010: c <= 9'b10111000;
				8'b1101101: c <= 9'b11111010;
				8'b100011: c <= 9'b10001100;
				8'b1110101: c <= 9'b1110000;
				8'b1111101: c <= 9'b100001011;
				8'b101001: c <= 9'b11111110;
				8'b1010010: c <= 9'b11000;
				8'b1011000: c <= 9'b11011101;
				8'b101110: c <= 9'b110000111;
				8'b1000001: c <= 9'b100100001;
				default: c <= 9'b0;
			endcase
			9'b101000100 : case(di)
				8'b1000011: c <= 9'b101;
				8'b101000: c <= 9'b10001000;
				8'b111010: c <= 9'b110000010;
				8'b110110: c <= 9'b111101100;
				8'b1100100: c <= 9'b101101000;
				8'b1000000: c <= 9'b10110110;
				8'b1110110: c <= 9'b101001100;
				8'b100101: c <= 9'b101110000;
				8'b101111: c <= 9'b110110101;
				8'b100110: c <= 9'b110100100;
				8'b1100011: c <= 9'b111100110;
				8'b1001000: c <= 9'b111110110;
				8'b111000: c <= 9'b100010011;
				8'b110001: c <= 9'b1000011;
				8'b1010111: c <= 9'b101001110;
				8'b1001110: c <= 9'b10111000;
				8'b1101010: c <= 9'b101110001;
				8'b1001001: c <= 9'b10100;
				8'b1100000: c <= 9'b10001101;
				8'b110111: c <= 9'b110101001;
				8'b1011101: c <= 9'b11111110;
				8'b1011011: c <= 9'b11010001;
				8'b111001: c <= 9'b1011001;
				8'b1001010: c <= 9'b100000011;
				8'b110011: c <= 9'b11100;
				8'b1101100: c <= 9'b101100111;
				8'b1110111: c <= 9'b111100100;
				8'b101011: c <= 9'b11100011;
				8'b1101011: c <= 9'b111011001;
				8'b111100: c <= 9'b1010001;
				8'b1000111: c <= 9'b10010101;
				8'b1011111: c <= 9'b100100101;
				8'b1110100: c <= 9'b110110100;
				8'b101101: c <= 9'b100110;
				8'b1010011: c <= 9'b1010000;
				8'b1100001: c <= 9'b111001100;
				8'b110101: c <= 9'b111100100;
				8'b1000100: c <= 9'b110011;
				8'b1010001: c <= 9'b11100101;
				8'b1010100: c <= 9'b11110011;
				8'b1100110: c <= 9'b100011101;
				8'b101010: c <= 9'b1100110;
				8'b1011110: c <= 9'b110001101;
				8'b1100111: c <= 9'b111001111;
				8'b1011010: c <= 9'b10110001;
				8'b1000010: c <= 9'b11011011;
				8'b111101: c <= 9'b110111111;
				8'b110000: c <= 9'b101000100;
				8'b111110: c <= 9'b10001100;
				8'b1100010: c <= 9'b11101;
				8'b1110000: c <= 9'b101000100;
				8'b1101001: c <= 9'b10100100;
				8'b1110011: c <= 9'b110111111;
				8'b1001100: c <= 9'b101000100;
				8'b100001: c <= 9'b10000110;
				8'b1000110: c <= 9'b110001000;
				8'b1110010: c <= 9'b111100101;
				8'b1010000: c <= 9'b110011000;
				8'b1111010: c <= 9'b1110111;
				8'b1010101: c <= 9'b10111011;
				8'b111011: c <= 9'b10000;
				8'b1001101: c <= 9'b10100100;
				8'b111111: c <= 9'b111100000;
				8'b1101110: c <= 9'b1011100;
				8'b1111011: c <= 9'b100011101;
				8'b1001011: c <= 9'b111100000;
				8'b1101111: c <= 9'b111110000;
				8'b1101000: c <= 9'b110011100;
				8'b101100: c <= 9'b101101110;
				8'b100100: c <= 9'b111011111;
				8'b1111000: c <= 9'b10111100;
				8'b1000101: c <= 9'b111111101;
				8'b1011001: c <= 9'b101100111;
				8'b110100: c <= 9'b110001101;
				8'b1111001: c <= 9'b1110001;
				8'b1110001: c <= 9'b1011000;
				8'b1001111: c <= 9'b111001100;
				8'b1100101: c <= 9'b10111001;
				8'b1111110: c <= 9'b1110101;
				8'b1111100: c <= 9'b110100110;
				8'b1010110: c <= 9'b10010;
				8'b110010: c <= 9'b1011011;
				8'b1101101: c <= 9'b1101000;
				8'b100011: c <= 9'b110110000;
				8'b1110101: c <= 9'b110000101;
				8'b1111101: c <= 9'b101010101;
				8'b101001: c <= 9'b101110111;
				8'b1010010: c <= 9'b1000100;
				8'b1011000: c <= 9'b101111111;
				8'b101110: c <= 9'b111101010;
				8'b1000001: c <= 9'b100010001;
				default: c <= 9'b0;
			endcase
			9'b111000111 : case(di)
				8'b1000011: c <= 9'b111000101;
				8'b101000: c <= 9'b110;
				8'b111010: c <= 9'b100111110;
				8'b110110: c <= 9'b11010011;
				8'b1100100: c <= 9'b101010100;
				8'b1000000: c <= 9'b100011010;
				8'b1110110: c <= 9'b100111011;
				8'b100101: c <= 9'b11111;
				8'b101111: c <= 9'b10111111;
				8'b100110: c <= 9'b110100111;
				8'b1100011: c <= 9'b110101111;
				8'b1001000: c <= 9'b111110101;
				8'b111000: c <= 9'b110011101;
				8'b110001: c <= 9'b110001000;
				8'b1010111: c <= 9'b10101;
				8'b1001110: c <= 9'b111010110;
				8'b1101010: c <= 9'b111100011;
				8'b1001001: c <= 9'b10110101;
				8'b1100000: c <= 9'b11000000;
				8'b110111: c <= 9'b1011100;
				8'b1011101: c <= 9'b110001110;
				8'b1011011: c <= 9'b101000101;
				8'b111001: c <= 9'b100010111;
				8'b1001010: c <= 9'b100110101;
				8'b110011: c <= 9'b1000100;
				8'b1101100: c <= 9'b11110001;
				8'b1110111: c <= 9'b100110000;
				8'b101011: c <= 9'b110111001;
				8'b1101011: c <= 9'b11100111;
				8'b111100: c <= 9'b10111001;
				8'b1000111: c <= 9'b1010111;
				8'b1011111: c <= 9'b11111010;
				8'b1110100: c <= 9'b1100001;
				8'b101101: c <= 9'b10111100;
				8'b1010011: c <= 9'b111000111;
				8'b1100001: c <= 9'b111001000;
				8'b110101: c <= 9'b1110010;
				8'b1000100: c <= 9'b110110010;
				8'b1010001: c <= 9'b10001111;
				8'b1010100: c <= 9'b111001001;
				8'b1100110: c <= 9'b111001110;
				8'b101010: c <= 9'b111100010;
				8'b1011110: c <= 9'b11000000;
				8'b1100111: c <= 9'b111000000;
				8'b1011010: c <= 9'b110000101;
				8'b1000010: c <= 9'b101;
				8'b111101: c <= 9'b10000011;
				8'b110000: c <= 9'b11010000;
				8'b111110: c <= 9'b100011111;
				8'b1100010: c <= 9'b1110100;
				8'b1110000: c <= 9'b100110101;
				8'b1101001: c <= 9'b1011010;
				8'b1110011: c <= 9'b100101010;
				8'b1001100: c <= 9'b100101100;
				8'b100001: c <= 9'b10011001;
				8'b1000110: c <= 9'b1000000;
				8'b1110010: c <= 9'b11101001;
				8'b1010000: c <= 9'b110111001;
				8'b1111010: c <= 9'b111101;
				8'b1010101: c <= 9'b110000010;
				8'b111011: c <= 9'b10010100;
				8'b1001101: c <= 9'b111;
				8'b111111: c <= 9'b10110100;
				8'b1101110: c <= 9'b101110111;
				8'b1111011: c <= 9'b11010010;
				8'b1001011: c <= 9'b100011010;
				8'b1101111: c <= 9'b100111100;
				8'b1101000: c <= 9'b100111011;
				8'b101100: c <= 9'b111101111;
				8'b100100: c <= 9'b100110100;
				8'b1111000: c <= 9'b100000111;
				8'b1000101: c <= 9'b100101000;
				8'b1011001: c <= 9'b1111101;
				8'b110100: c <= 9'b100101110;
				8'b1111001: c <= 9'b10110010;
				8'b1110001: c <= 9'b100100;
				8'b1001111: c <= 9'b100110000;
				8'b1100101: c <= 9'b10010011;
				8'b1111110: c <= 9'b1010001;
				8'b1111100: c <= 9'b110011101;
				8'b1010110: c <= 9'b10011011;
				8'b110010: c <= 9'b110101001;
				8'b1101101: c <= 9'b101010010;
				8'b100011: c <= 9'b100001111;
				8'b1110101: c <= 9'b11100;
				8'b1111101: c <= 9'b101011111;
				8'b101001: c <= 9'b110000010;
				8'b1010010: c <= 9'b100000010;
				8'b1011000: c <= 9'b100100110;
				8'b101110: c <= 9'b11011010;
				8'b1000001: c <= 9'b1111101;
				default: c <= 9'b0;
			endcase
			9'b111010110 : case(di)
				8'b1000011: c <= 9'b101001000;
				8'b101000: c <= 9'b1101101;
				8'b111010: c <= 9'b101100;
				8'b110110: c <= 9'b1100001;
				8'b1100100: c <= 9'b10000000;
				8'b1000000: c <= 9'b100111110;
				8'b1110110: c <= 9'b101101000;
				8'b100101: c <= 9'b110101001;
				8'b101111: c <= 9'b10100011;
				8'b100110: c <= 9'b100110011;
				8'b1100011: c <= 9'b10010100;
				8'b1001000: c <= 9'b100001101;
				8'b111000: c <= 9'b101001;
				8'b110001: c <= 9'b110000111;
				8'b1010111: c <= 9'b100110100;
				8'b1001110: c <= 9'b111000101;
				8'b1101010: c <= 9'b10000011;
				8'b1001001: c <= 9'b10101110;
				8'b1100000: c <= 9'b100011111;
				8'b110111: c <= 9'b11100111;
				8'b1011101: c <= 9'b11001000;
				8'b1011011: c <= 9'b10010111;
				8'b111001: c <= 9'b10111010;
				8'b1001010: c <= 9'b10110101;
				8'b110011: c <= 9'b100001001;
				8'b1101100: c <= 9'b100111110;
				8'b1110111: c <= 9'b1010001;
				8'b101011: c <= 9'b101111110;
				8'b1101011: c <= 9'b110100101;
				8'b111100: c <= 9'b11000011;
				8'b1000111: c <= 9'b10010011;
				8'b1011111: c <= 9'b100000011;
				8'b1110100: c <= 9'b11100010;
				8'b101101: c <= 9'b101010100;
				8'b1010011: c <= 9'b101101010;
				8'b1100001: c <= 9'b11101;
				8'b110101: c <= 9'b110100010;
				8'b1000100: c <= 9'b101010010;
				8'b1010001: c <= 9'b111100000;
				8'b1010100: c <= 9'b101000011;
				8'b1100110: c <= 9'b110100110;
				8'b101010: c <= 9'b10110010;
				8'b1011110: c <= 9'b11000001;
				8'b1100111: c <= 9'b101011111;
				8'b1011010: c <= 9'b111011;
				8'b1000010: c <= 9'b100011101;
				8'b111101: c <= 9'b101101001;
				8'b110000: c <= 9'b101101100;
				8'b111110: c <= 9'b10100101;
				8'b1100010: c <= 9'b1111111;
				8'b1110000: c <= 9'b101011101;
				8'b1101001: c <= 9'b11111010;
				8'b1110011: c <= 9'b101000;
				8'b1001100: c <= 9'b110000110;
				8'b100001: c <= 9'b10101101;
				8'b1000110: c <= 9'b111001101;
				8'b1110010: c <= 9'b10101001;
				8'b1010000: c <= 9'b1101001;
				8'b1111010: c <= 9'b10001001;
				8'b1010101: c <= 9'b10010110;
				8'b111011: c <= 9'b101100010;
				8'b1001101: c <= 9'b100000101;
				8'b111111: c <= 9'b11101101;
				8'b1101110: c <= 9'b10101110;
				8'b1111011: c <= 9'b11110110;
				8'b1001011: c <= 9'b100011011;
				8'b1101111: c <= 9'b100000100;
				8'b1101000: c <= 9'b11100010;
				8'b101100: c <= 9'b11011101;
				8'b100100: c <= 9'b111100011;
				8'b1111000: c <= 9'b100011000;
				8'b1000101: c <= 9'b1111010;
				8'b1011001: c <= 9'b100100001;
				8'b110100: c <= 9'b10101011;
				8'b1111001: c <= 9'b11000110;
				8'b1110001: c <= 9'b101100110;
				8'b1001111: c <= 9'b10110;
				8'b1100101: c <= 9'b11101;
				8'b1111110: c <= 9'b11111011;
				8'b1111100: c <= 9'b101000111;
				8'b1010110: c <= 9'b111101;
				8'b110010: c <= 9'b110000010;
				8'b1101101: c <= 9'b111101001;
				8'b100011: c <= 9'b110001110;
				8'b1110101: c <= 9'b100101101;
				8'b1111101: c <= 9'b111100;
				8'b101001: c <= 9'b11110011;
				8'b1010010: c <= 9'b1110100;
				8'b1011000: c <= 9'b1001001;
				8'b101110: c <= 9'b1110101;
				8'b1000001: c <= 9'b111101001;
				default: c <= 9'b0;
			endcase
			9'b100101001 : case(di)
				8'b1000011: c <= 9'b100010110;
				8'b101000: c <= 9'b101010010;
				8'b111010: c <= 9'b100100101;
				8'b110110: c <= 9'b111001001;
				8'b1100100: c <= 9'b110100100;
				8'b1000000: c <= 9'b10001010;
				8'b1110110: c <= 9'b111000100;
				8'b100101: c <= 9'b11110111;
				8'b101111: c <= 9'b100100110;
				8'b100110: c <= 9'b110110100;
				8'b1100011: c <= 9'b1001000;
				8'b1001000: c <= 9'b101010001;
				8'b111000: c <= 9'b10010101;
				8'b110001: c <= 9'b101101000;
				8'b1010111: c <= 9'b111010111;
				8'b1001110: c <= 9'b111100111;
				8'b1101010: c <= 9'b1110000;
				8'b1001001: c <= 9'b10011100;
				8'b1100000: c <= 9'b11111000;
				8'b110111: c <= 9'b11100011;
				8'b1011101: c <= 9'b10111110;
				8'b1011011: c <= 9'b101111111;
				8'b111001: c <= 9'b100000010;
				8'b1001010: c <= 9'b11000111;
				8'b110011: c <= 9'b100000101;
				8'b1101100: c <= 9'b11010101;
				8'b1110111: c <= 9'b10111011;
				8'b101011: c <= 9'b100000110;
				8'b1101011: c <= 9'b110110100;
				8'b111100: c <= 9'b110011000;
				8'b1000111: c <= 9'b101010110;
				8'b1011111: c <= 9'b100101010;
				8'b1110100: c <= 9'b100010000;
				8'b101101: c <= 9'b100010100;
				8'b1010011: c <= 9'b1111100;
				8'b1100001: c <= 9'b111001110;
				8'b110101: c <= 9'b100100010;
				8'b1000100: c <= 9'b111001111;
				8'b1010001: c <= 9'b111100;
				8'b1010100: c <= 9'b111010001;
				8'b1100110: c <= 9'b100010101;
				8'b101010: c <= 9'b10111;
				8'b1011110: c <= 9'b1000100;
				8'b1100111: c <= 9'b1001111;
				8'b1011010: c <= 9'b1001100;
				8'b1000010: c <= 9'b1010011;
				8'b111101: c <= 9'b111;
				8'b110000: c <= 9'b11111001;
				8'b111110: c <= 9'b11011011;
				8'b1100010: c <= 9'b101011110;
				8'b1110000: c <= 9'b100110011;
				8'b1101001: c <= 9'b1010000;
				8'b1110011: c <= 9'b11000011;
				8'b1001100: c <= 9'b101101011;
				8'b100001: c <= 9'b10011010;
				8'b1000110: c <= 9'b1101001;
				8'b1110010: c <= 9'b10011111;
				8'b1010000: c <= 9'b1111101;
				8'b1111010: c <= 9'b10001111;
				8'b1010101: c <= 9'b111100;
				8'b111011: c <= 9'b110000000;
				8'b1001101: c <= 9'b110110000;
				8'b111111: c <= 9'b110101011;
				8'b1101110: c <= 9'b11000;
				8'b1111011: c <= 9'b110100100;
				8'b1001011: c <= 9'b111101;
				8'b1101111: c <= 9'b1011111;
				8'b1101000: c <= 9'b11110001;
				8'b101100: c <= 9'b100110010;
				8'b100100: c <= 9'b111111110;
				8'b1111000: c <= 9'b10010000;
				8'b1000101: c <= 9'b100101111;
				8'b1011001: c <= 9'b111111111;
				8'b110100: c <= 9'b100100;
				8'b1111001: c <= 9'b11111100;
				8'b1110001: c <= 9'b101011000;
				8'b1001111: c <= 9'b1110000;
				8'b1100101: c <= 9'b11010;
				8'b1111110: c <= 9'b10011101;
				8'b1111100: c <= 9'b11110000;
				8'b1010110: c <= 9'b10100110;
				8'b110010: c <= 9'b11001;
				8'b1101101: c <= 9'b101011001;
				8'b100011: c <= 9'b110000101;
				8'b1110101: c <= 9'b100011011;
				8'b1111101: c <= 9'b110011010;
				8'b101001: c <= 9'b10000110;
				8'b1010010: c <= 9'b110111001;
				8'b1011000: c <= 9'b101000011;
				8'b101110: c <= 9'b100000010;
				8'b1000001: c <= 9'b111000;
				default: c <= 9'b0;
			endcase
			9'b1001101 : case(di)
				8'b1000011: c <= 9'b100011000;
				8'b101000: c <= 9'b110110;
				8'b111010: c <= 9'b100111000;
				8'b110110: c <= 9'b111111;
				8'b1100100: c <= 9'b10111110;
				8'b1000000: c <= 9'b111111110;
				8'b1110110: c <= 9'b1011000;
				8'b100101: c <= 9'b111010000;
				8'b101111: c <= 9'b110011011;
				8'b100110: c <= 9'b101110100;
				8'b1100011: c <= 9'b1110111;
				8'b1001000: c <= 9'b111111111;
				8'b111000: c <= 9'b101011010;
				8'b110001: c <= 9'b110001111;
				8'b1010111: c <= 9'b100110011;
				8'b1001110: c <= 9'b110000010;
				8'b1101010: c <= 9'b10010110;
				8'b1001001: c <= 9'b101100100;
				8'b1100000: c <= 9'b111001110;
				8'b110111: c <= 9'b111000100;
				8'b1011101: c <= 9'b100010011;
				8'b1011011: c <= 9'b10010001;
				8'b111001: c <= 9'b101100011;
				8'b1001010: c <= 9'b100100101;
				8'b110011: c <= 9'b10111;
				8'b1101100: c <= 9'b101001001;
				8'b1110111: c <= 9'b1010000;
				8'b101011: c <= 9'b110000000;
				8'b1101011: c <= 9'b10011011;
				8'b111100: c <= 9'b111100001;
				8'b1000111: c <= 9'b101011111;
				8'b1011111: c <= 9'b101101110;
				8'b1110100: c <= 9'b110011100;
				8'b101101: c <= 9'b101110011;
				8'b1010011: c <= 9'b111100010;
				8'b1100001: c <= 9'b110101110;
				8'b110101: c <= 9'b110001110;
				8'b1000100: c <= 9'b100010111;
				8'b1010001: c <= 9'b101110101;
				8'b1010100: c <= 9'b101110000;
				8'b1100110: c <= 9'b110010111;
				8'b101010: c <= 9'b10000101;
				8'b1011110: c <= 9'b10110111;
				8'b1100111: c <= 9'b100110;
				8'b1011010: c <= 9'b111101110;
				8'b1000010: c <= 9'b10100011;
				8'b111101: c <= 9'b11001;
				8'b110000: c <= 9'b10011011;
				8'b111110: c <= 9'b1101110;
				8'b1100010: c <= 9'b1001011;
				8'b1110000: c <= 9'b10110011;
				8'b1101001: c <= 9'b111111110;
				8'b1110011: c <= 9'b101110011;
				8'b1001100: c <= 9'b110110000;
				8'b100001: c <= 9'b1111000;
				8'b1000110: c <= 9'b100110;
				8'b1110010: c <= 9'b11111011;
				8'b1010000: c <= 9'b110101101;
				8'b1111010: c <= 9'b110100010;
				8'b1010101: c <= 9'b1101;
				8'b111011: c <= 9'b111110000;
				8'b1001101: c <= 9'b111011010;
				8'b111111: c <= 9'b1101000;
				8'b1101110: c <= 9'b100101000;
				8'b1111011: c <= 9'b110;
				8'b1001011: c <= 9'b100111;
				8'b1101111: c <= 9'b10101011;
				8'b1101000: c <= 9'b100001111;
				8'b101100: c <= 9'b1001010;
				8'b100100: c <= 9'b11010111;
				8'b1111000: c <= 9'b100010;
				8'b1000101: c <= 9'b100111011;
				8'b1011001: c <= 9'b101111111;
				8'b110100: c <= 9'b101001;
				8'b1111001: c <= 9'b10110101;
				8'b1110001: c <= 9'b10010101;
				8'b1001111: c <= 9'b101011;
				8'b1100101: c <= 9'b100010;
				8'b1111110: c <= 9'b10100110;
				8'b1111100: c <= 9'b10000110;
				8'b1010110: c <= 9'b101100000;
				8'b110010: c <= 9'b100011101;
				8'b1101101: c <= 9'b110100111;
				8'b100011: c <= 9'b110110011;
				8'b1110101: c <= 9'b1010001;
				8'b1111101: c <= 9'b10111001;
				8'b101001: c <= 9'b1010000;
				8'b1010010: c <= 9'b100001101;
				8'b1011000: c <= 9'b11001100;
				8'b101110: c <= 9'b100101110;
				8'b1000001: c <= 9'b10111011;
				default: c <= 9'b0;
			endcase
			9'b101000110 : case(di)
				8'b1000011: c <= 9'b111000011;
				8'b101000: c <= 9'b100100011;
				8'b111010: c <= 9'b111000100;
				8'b110110: c <= 9'b100000111;
				8'b1100100: c <= 9'b110100101;
				8'b1000000: c <= 9'b101100010;
				8'b1110110: c <= 9'b101001001;
				8'b100101: c <= 9'b101001110;
				8'b101111: c <= 9'b1100011;
				8'b100110: c <= 9'b101001110;
				8'b1100011: c <= 9'b1011010;
				8'b1001000: c <= 9'b11100101;
				8'b111000: c <= 9'b11001111;
				8'b110001: c <= 9'b100000000;
				8'b1010111: c <= 9'b100000001;
				8'b1001110: c <= 9'b10100000;
				8'b1101010: c <= 9'b11111001;
				8'b1001001: c <= 9'b111001100;
				8'b1100000: c <= 9'b11101;
				8'b110111: c <= 9'b101101000;
				8'b1011101: c <= 9'b110101010;
				8'b1011011: c <= 9'b11001001;
				8'b111001: c <= 9'b1111001;
				8'b1001010: c <= 9'b100000111;
				8'b110011: c <= 9'b101001010;
				8'b1101100: c <= 9'b110101101;
				8'b1110111: c <= 9'b100111100;
				8'b101011: c <= 9'b11001;
				8'b1101011: c <= 9'b100110;
				8'b111100: c <= 9'b111100100;
				8'b1000111: c <= 9'b10101100;
				8'b1011111: c <= 9'b100001011;
				8'b1110100: c <= 9'b111000010;
				8'b101101: c <= 9'b10110100;
				8'b1010011: c <= 9'b101010001;
				8'b1100001: c <= 9'b110011111;
				8'b110101: c <= 9'b101010000;
				8'b1000100: c <= 9'b1111000;
				8'b1010001: c <= 9'b110011011;
				8'b1010100: c <= 9'b100110;
				8'b1100110: c <= 9'b111010010;
				8'b101010: c <= 9'b111001001;
				8'b1011110: c <= 9'b111100110;
				8'b1100111: c <= 9'b100111010;
				8'b1011010: c <= 9'b1111111;
				8'b1000010: c <= 9'b100010100;
				8'b111101: c <= 9'b111100000;
				8'b110000: c <= 9'b101010110;
				8'b111110: c <= 9'b10000011;
				8'b1100010: c <= 9'b11110111;
				8'b1110000: c <= 9'b11110000;
				8'b1101001: c <= 9'b101010100;
				8'b1110011: c <= 9'b1110100;
				8'b1001100: c <= 9'b100100000;
				8'b100001: c <= 9'b101011011;
				8'b1000110: c <= 9'b101001010;
				8'b1110010: c <= 9'b101010101;
				8'b1010000: c <= 9'b100000011;
				8'b1111010: c <= 9'b101110000;
				8'b1010101: c <= 9'b100001001;
				8'b111011: c <= 9'b11001101;
				8'b1001101: c <= 9'b10000001;
				8'b111111: c <= 9'b1111010;
				8'b1101110: c <= 9'b10011000;
				8'b1111011: c <= 9'b10101100;
				8'b1001011: c <= 9'b11110011;
				8'b1101111: c <= 9'b10110001;
				8'b1101000: c <= 9'b1101111;
				8'b101100: c <= 9'b101111000;
				8'b100100: c <= 9'b100011100;
				8'b1111000: c <= 9'b1101000;
				8'b1000101: c <= 9'b10100010;
				8'b1011001: c <= 9'b1100001;
				8'b110100: c <= 9'b10100101;
				8'b1111001: c <= 9'b100101110;
				8'b1110001: c <= 9'b10100110;
				8'b1001111: c <= 9'b101001100;
				8'b1100101: c <= 9'b11100101;
				8'b1111110: c <= 9'b100000000;
				8'b1111100: c <= 9'b100010101;
				8'b1010110: c <= 9'b111111010;
				8'b110010: c <= 9'b110011111;
				8'b1101101: c <= 9'b110010;
				8'b100011: c <= 9'b110010011;
				8'b1110101: c <= 9'b100011001;
				8'b1111101: c <= 9'b101101010;
				8'b101001: c <= 9'b1001011;
				8'b1010010: c <= 9'b110001011;
				8'b1011000: c <= 9'b100010000;
				8'b101110: c <= 9'b110111000;
				8'b1000001: c <= 9'b100001110;
				default: c <= 9'b0;
			endcase
			9'b1011000 : case(di)
				8'b1000011: c <= 9'b10100101;
				8'b101000: c <= 9'b101110001;
				8'b111010: c <= 9'b111111101;
				8'b110110: c <= 9'b101101011;
				8'b1100100: c <= 9'b1000100;
				8'b1000000: c <= 9'b101011001;
				8'b1110110: c <= 9'b1100100;
				8'b100101: c <= 9'b100011101;
				8'b101111: c <= 9'b111110101;
				8'b100110: c <= 9'b100101001;
				8'b1100011: c <= 9'b10011001;
				8'b1001000: c <= 9'b111100110;
				8'b111000: c <= 9'b100110101;
				8'b110001: c <= 9'b111100000;
				8'b1010111: c <= 9'b11001101;
				8'b1001110: c <= 9'b1101110;
				8'b1101010: c <= 9'b11100000;
				8'b1001001: c <= 9'b100001100;
				8'b1100000: c <= 9'b111000;
				8'b110111: c <= 9'b10011111;
				8'b1011101: c <= 9'b11011001;
				8'b1011011: c <= 9'b110110110;
				8'b111001: c <= 9'b1100001;
				8'b1001010: c <= 9'b100110011;
				8'b110011: c <= 9'b1000011;
				8'b1101100: c <= 9'b100010100;
				8'b1110111: c <= 9'b1000010;
				8'b101011: c <= 9'b101100;
				8'b1101011: c <= 9'b11010000;
				8'b111100: c <= 9'b111001;
				8'b1000111: c <= 9'b110000111;
				8'b1011111: c <= 9'b111101101;
				8'b1110100: c <= 9'b10100010;
				8'b101101: c <= 9'b1010000;
				8'b1010011: c <= 9'b110001101;
				8'b1100001: c <= 9'b101010001;
				8'b110101: c <= 9'b11001001;
				8'b1000100: c <= 9'b101010001;
				8'b1010001: c <= 9'b100111011;
				8'b1010100: c <= 9'b10000010;
				8'b1100110: c <= 9'b101101110;
				8'b101010: c <= 9'b1000001;
				8'b1011110: c <= 9'b101000110;
				8'b1100111: c <= 9'b1011000;
				8'b1011010: c <= 9'b10101001;
				8'b1000010: c <= 9'b111111001;
				8'b111101: c <= 9'b10100000;
				8'b110000: c <= 9'b1101101;
				8'b111110: c <= 9'b100000111;
				8'b1100010: c <= 9'b111111110;
				8'b1110000: c <= 9'b10101100;
				8'b1101001: c <= 9'b111001111;
				8'b1110011: c <= 9'b110010100;
				8'b1001100: c <= 9'b110100001;
				8'b100001: c <= 9'b110011010;
				8'b1000110: c <= 9'b1011011;
				8'b1110010: c <= 9'b110110011;
				8'b1010000: c <= 9'b101010010;
				8'b1111010: c <= 9'b110111111;
				8'b1010101: c <= 9'b10100011;
				8'b111011: c <= 9'b110100;
				8'b1001101: c <= 9'b10100110;
				8'b111111: c <= 9'b101101011;
				8'b1101110: c <= 9'b110100101;
				8'b1111011: c <= 9'b1100000;
				8'b1001011: c <= 9'b100101001;
				8'b1101111: c <= 9'b111110101;
				8'b1101000: c <= 9'b100110011;
				8'b101100: c <= 9'b110010001;
				8'b100100: c <= 9'b111101010;
				8'b1111000: c <= 9'b101100011;
				8'b1000101: c <= 9'b10000110;
				8'b1011001: c <= 9'b1101111;
				8'b110100: c <= 9'b1000011;
				8'b1111001: c <= 9'b10110;
				8'b1110001: c <= 9'b111101101;
				8'b1001111: c <= 9'b100101110;
				8'b1100101: c <= 9'b1001101;
				8'b1111110: c <= 9'b110001001;
				8'b1111100: c <= 9'b11100110;
				8'b1010110: c <= 9'b110000011;
				8'b110010: c <= 9'b10000000;
				8'b1101101: c <= 9'b100011011;
				8'b100011: c <= 9'b111110000;
				8'b1110101: c <= 9'b110010001;
				8'b1111101: c <= 9'b111001100;
				8'b101001: c <= 9'b111000110;
				8'b1010010: c <= 9'b1011001;
				8'b1011000: c <= 9'b10110111;
				8'b101110: c <= 9'b10101001;
				8'b1000001: c <= 9'b1001001;
				default: c <= 9'b0;
			endcase
			9'b11110101 : case(di)
				8'b1000011: c <= 9'b100110100;
				8'b101000: c <= 9'b111101010;
				8'b111010: c <= 9'b10010100;
				8'b110110: c <= 9'b100001111;
				8'b1100100: c <= 9'b101101010;
				8'b1000000: c <= 9'b11000011;
				8'b1110110: c <= 9'b100011;
				8'b100101: c <= 9'b100111111;
				8'b101111: c <= 9'b11000001;
				8'b100110: c <= 9'b111111010;
				8'b1100011: c <= 9'b11100011;
				8'b1001000: c <= 9'b111110011;
				8'b111000: c <= 9'b1000011;
				8'b110001: c <= 9'b101011000;
				8'b1010111: c <= 9'b101001111;
				8'b1001110: c <= 9'b100101100;
				8'b1101010: c <= 9'b10000011;
				8'b1001001: c <= 9'b101001100;
				8'b1100000: c <= 9'b1000100;
				8'b110111: c <= 9'b111100110;
				8'b1011101: c <= 9'b100001010;
				8'b1011011: c <= 9'b11111100;
				8'b111001: c <= 9'b1100001;
				8'b1001010: c <= 9'b11010100;
				8'b110011: c <= 9'b100011011;
				8'b1101100: c <= 9'b11010011;
				8'b1110111: c <= 9'b110101001;
				8'b101011: c <= 9'b10010;
				8'b1101011: c <= 9'b101101010;
				8'b111100: c <= 9'b101001110;
				8'b1000111: c <= 9'b110010110;
				8'b1011111: c <= 9'b11101111;
				8'b1110100: c <= 9'b10101000;
				8'b101101: c <= 9'b1011010;
				8'b1010011: c <= 9'b100110011;
				8'b1100001: c <= 9'b111101100;
				8'b110101: c <= 9'b11111010;
				8'b1000100: c <= 9'b110110;
				8'b1010001: c <= 9'b110100111;
				8'b1010100: c <= 9'b111111000;
				8'b1100110: c <= 9'b10100010;
				8'b101010: c <= 9'b100010101;
				8'b1011110: c <= 9'b1101111;
				8'b1100111: c <= 9'b11000111;
				8'b1011010: c <= 9'b110001011;
				8'b1000010: c <= 9'b100010110;
				8'b111101: c <= 9'b110110;
				8'b110000: c <= 9'b11101101;
				8'b111110: c <= 9'b100011010;
				8'b1100010: c <= 9'b101110111;
				8'b1110000: c <= 9'b10110;
				8'b1101001: c <= 9'b101100000;
				8'b1110011: c <= 9'b1000010;
				8'b1001100: c <= 9'b11100000;
				8'b100001: c <= 9'b111010111;
				8'b1000110: c <= 9'b100110;
				8'b1110010: c <= 9'b10011111;
				8'b1010000: c <= 9'b1000001;
				8'b1111010: c <= 9'b11110100;
				8'b1010101: c <= 9'b110001001;
				8'b111011: c <= 9'b1110000;
				8'b1001101: c <= 9'b10100000;
				8'b111111: c <= 9'b101010100;
				8'b1101110: c <= 9'b101101100;
				8'b1111011: c <= 9'b110000011;
				8'b1001011: c <= 9'b10010110;
				8'b1101111: c <= 9'b111101001;
				8'b1101000: c <= 9'b11101001;
				8'b101100: c <= 9'b1110111;
				8'b100100: c <= 9'b111100110;
				8'b1111000: c <= 9'b11110100;
				8'b1000101: c <= 9'b111001010;
				8'b1011001: c <= 9'b11000001;
				8'b110100: c <= 9'b10000101;
				8'b1111001: c <= 9'b100100101;
				8'b1110001: c <= 9'b101100110;
				8'b1001111: c <= 9'b100111101;
				8'b1100101: c <= 9'b100001100;
				8'b1111110: c <= 9'b110010001;
				8'b1111100: c <= 9'b101000110;
				8'b1010110: c <= 9'b100100011;
				8'b110010: c <= 9'b111000011;
				8'b1101101: c <= 9'b100001101;
				8'b100011: c <= 9'b111100010;
				8'b1110101: c <= 9'b111000100;
				8'b1111101: c <= 9'b111010000;
				8'b101001: c <= 9'b11001011;
				8'b1010010: c <= 9'b110110100;
				8'b1011000: c <= 9'b11001;
				8'b101110: c <= 9'b1110011;
				8'b1000001: c <= 9'b10;
				default: c <= 9'b0;
			endcase
			9'b1010000 : case(di)
				8'b1000011: c <= 9'b10001000;
				8'b101000: c <= 9'b110100101;
				8'b111010: c <= 9'b101101101;
				8'b110110: c <= 9'b101010001;
				8'b1100100: c <= 9'b11100010;
				8'b1000000: c <= 9'b111100000;
				8'b1110110: c <= 9'b10010111;
				8'b100101: c <= 9'b111000110;
				8'b101111: c <= 9'b101101;
				8'b100110: c <= 9'b111001110;
				8'b1100011: c <= 9'b1000;
				8'b1001000: c <= 9'b1011100;
				8'b111000: c <= 9'b101101;
				8'b110001: c <= 9'b10000011;
				8'b1010111: c <= 9'b101110000;
				8'b1001110: c <= 9'b111111001;
				8'b1101010: c <= 9'b101010110;
				8'b1001001: c <= 9'b101010001;
				8'b1100000: c <= 9'b101010111;
				8'b110111: c <= 9'b101000111;
				8'b1011101: c <= 9'b100101011;
				8'b1011011: c <= 9'b1111000;
				8'b111001: c <= 9'b111111010;
				8'b1001010: c <= 9'b111010;
				8'b110011: c <= 9'b1001100;
				8'b1101100: c <= 9'b111010001;
				8'b1110111: c <= 9'b10010110;
				8'b101011: c <= 9'b11000111;
				8'b1101011: c <= 9'b110001010;
				8'b111100: c <= 9'b101000001;
				8'b1000111: c <= 9'b111011011;
				8'b1011111: c <= 9'b100110010;
				8'b1110100: c <= 9'b11111110;
				8'b101101: c <= 9'b111111001;
				8'b1010011: c <= 9'b11011001;
				8'b1100001: c <= 9'b100011101;
				8'b110101: c <= 9'b110101;
				8'b1000100: c <= 9'b1110101;
				8'b1010001: c <= 9'b101001110;
				8'b1010100: c <= 9'b10111111;
				8'b1100110: c <= 9'b1011110;
				8'b101010: c <= 9'b100111101;
				8'b1011110: c <= 9'b11001101;
				8'b1100111: c <= 9'b11001010;
				8'b1011010: c <= 9'b11010000;
				8'b1000010: c <= 9'b110000011;
				8'b111101: c <= 9'b101100011;
				8'b110000: c <= 9'b11010100;
				8'b111110: c <= 9'b11011100;
				8'b1100010: c <= 9'b110101001;
				8'b1110000: c <= 9'b101001;
				8'b1101001: c <= 9'b100100101;
				8'b1110011: c <= 9'b101000001;
				8'b1001100: c <= 9'b111111;
				8'b100001: c <= 9'b110001011;
				8'b1000110: c <= 9'b11010010;
				8'b1110010: c <= 9'b101010000;
				8'b1010000: c <= 9'b101111110;
				8'b1111010: c <= 9'b100101000;
				8'b1010101: c <= 9'b11001110;
				8'b111011: c <= 9'b110101111;
				8'b1001101: c <= 9'b10010001;
				8'b111111: c <= 9'b1111010;
				8'b1101110: c <= 9'b10011101;
				8'b1111011: c <= 9'b101000010;
				8'b1001011: c <= 9'b1110111;
				8'b1101111: c <= 9'b100111111;
				8'b1101000: c <= 9'b101101010;
				8'b101100: c <= 9'b111001110;
				8'b100100: c <= 9'b111000011;
				8'b1111000: c <= 9'b100011100;
				8'b1000101: c <= 9'b101011010;
				8'b1011001: c <= 9'b110000000;
				8'b110100: c <= 9'b10101000;
				8'b1111001: c <= 9'b101001100;
				8'b1110001: c <= 9'b11100100;
				8'b1001111: c <= 9'b1011110;
				8'b1100101: c <= 9'b110001100;
				8'b1111110: c <= 9'b1001100;
				8'b1111100: c <= 9'b1100101;
				8'b1010110: c <= 9'b111101000;
				8'b110010: c <= 9'b11000100;
				8'b1101101: c <= 9'b100000111;
				8'b100011: c <= 9'b10000111;
				8'b1110101: c <= 9'b111111011;
				8'b1111101: c <= 9'b110010010;
				8'b101001: c <= 9'b11100101;
				8'b1010010: c <= 9'b111101001;
				8'b1011000: c <= 9'b100100000;
				8'b101110: c <= 9'b101011101;
				8'b1000001: c <= 9'b110010;
				default: c <= 9'b0;
			endcase
			9'b101100 : case(di)
				8'b1000011: c <= 9'b100101;
				8'b101000: c <= 9'b1101000;
				8'b111010: c <= 9'b1001110;
				8'b110110: c <= 9'b101001011;
				8'b1100100: c <= 9'b100101100;
				8'b1000000: c <= 9'b11001;
				8'b1110110: c <= 9'b111110011;
				8'b100101: c <= 9'b1100;
				8'b101111: c <= 9'b1100010;
				8'b100110: c <= 9'b100000010;
				8'b1100011: c <= 9'b100011001;
				8'b1001000: c <= 9'b1101010;
				8'b111000: c <= 9'b11001100;
				8'b110001: c <= 9'b1100101;
				8'b1010111: c <= 9'b101010110;
				8'b1001110: c <= 9'b10110;
				8'b1101010: c <= 9'b110101101;
				8'b1001001: c <= 9'b1000000;
				8'b1100000: c <= 9'b110010101;
				8'b110111: c <= 9'b10111;
				8'b1011101: c <= 9'b111000100;
				8'b1011011: c <= 9'b11010111;
				8'b111001: c <= 9'b111110110;
				8'b1001010: c <= 9'b10000000;
				8'b110011: c <= 9'b1001111;
				8'b1101100: c <= 9'b101010110;
				8'b1110111: c <= 9'b110011010;
				8'b101011: c <= 9'b101101100;
				8'b1101011: c <= 9'b11000110;
				8'b111100: c <= 9'b11001101;
				8'b1000111: c <= 9'b11110;
				8'b1011111: c <= 9'b11101101;
				8'b1110100: c <= 9'b100011011;
				8'b101101: c <= 9'b11011101;
				8'b1010011: c <= 9'b100111110;
				8'b1100001: c <= 9'b111100000;
				8'b110101: c <= 9'b110010110;
				8'b1000100: c <= 9'b1100011;
				8'b1010001: c <= 9'b110100100;
				8'b1010100: c <= 9'b100100001;
				8'b1100110: c <= 9'b110001111;
				8'b101010: c <= 9'b111111111;
				8'b1011110: c <= 9'b100001101;
				8'b1100111: c <= 9'b111100000;
				8'b1011010: c <= 9'b110000011;
				8'b1000010: c <= 9'b101010110;
				8'b111101: c <= 9'b100100;
				8'b110000: c <= 9'b110011001;
				8'b111110: c <= 9'b101100000;
				8'b1100010: c <= 9'b110111111;
				8'b1110000: c <= 9'b1000001;
				8'b1101001: c <= 9'b11110101;
				8'b1110011: c <= 9'b111011110;
				8'b1001100: c <= 9'b10111010;
				8'b100001: c <= 9'b1001001;
				8'b1000110: c <= 9'b110111110;
				8'b1110010: c <= 9'b101000110;
				8'b1010000: c <= 9'b111100000;
				8'b1111010: c <= 9'b11111010;
				8'b1010101: c <= 9'b110010100;
				8'b111011: c <= 9'b110001011;
				8'b1001101: c <= 9'b1001011;
				8'b111111: c <= 9'b1110111;
				8'b1101110: c <= 9'b100101000;
				8'b1111011: c <= 9'b111110011;
				8'b1001011: c <= 9'b110100101;
				8'b1101111: c <= 9'b110001010;
				8'b1101000: c <= 9'b101101111;
				8'b101100: c <= 9'b1000100;
				8'b100100: c <= 9'b110001101;
				8'b1111000: c <= 9'b111111;
				8'b1000101: c <= 9'b1010000;
				8'b1011001: c <= 9'b100010001;
				8'b110100: c <= 9'b101100101;
				8'b1111001: c <= 9'b111000000;
				8'b1110001: c <= 9'b100110110;
				8'b1001111: c <= 9'b10100010;
				8'b1100101: c <= 9'b100001101;
				8'b1111110: c <= 9'b11;
				8'b1111100: c <= 9'b10100011;
				8'b1010110: c <= 9'b101101000;
				8'b110010: c <= 9'b10001011;
				8'b1101101: c <= 9'b101011010;
				8'b100011: c <= 9'b10011;
				8'b1110101: c <= 9'b111111011;
				8'b1111101: c <= 9'b101011011;
				8'b101001: c <= 9'b10100;
				8'b1010010: c <= 9'b110011010;
				8'b1011000: c <= 9'b11011011;
				8'b101110: c <= 9'b100111100;
				8'b1000001: c <= 9'b11000011;
				default: c <= 9'b0;
			endcase
			9'b11001010 : case(di)
				8'b1000011: c <= 9'b10111010;
				8'b101000: c <= 9'b10010011;
				8'b111010: c <= 9'b11011110;
				8'b110110: c <= 9'b110010100;
				8'b1100100: c <= 9'b10010011;
				8'b1000000: c <= 9'b11011110;
				8'b1110110: c <= 9'b111101000;
				8'b100101: c <= 9'b10001011;
				8'b101111: c <= 9'b100001010;
				8'b100110: c <= 9'b101000010;
				8'b1100011: c <= 9'b111000;
				8'b1001000: c <= 9'b11111101;
				8'b111000: c <= 9'b1;
				8'b110001: c <= 9'b10000111;
				8'b1010111: c <= 9'b100011001;
				8'b1001110: c <= 9'b100001001;
				8'b1101010: c <= 9'b100011;
				8'b1001001: c <= 9'b101011110;
				8'b1100000: c <= 9'b110110111;
				8'b110111: c <= 9'b101011110;
				8'b1011101: c <= 9'b11011010;
				8'b1011011: c <= 9'b101111001;
				8'b111001: c <= 9'b10001111;
				8'b1001010: c <= 9'b10100;
				8'b110011: c <= 9'b111110110;
				8'b1101100: c <= 9'b110011101;
				8'b1110111: c <= 9'b111010010;
				8'b101011: c <= 9'b110011001;
				8'b1101011: c <= 9'b10101;
				8'b111100: c <= 9'b101101100;
				8'b1000111: c <= 9'b1;
				8'b1011111: c <= 9'b100110100;
				8'b1110100: c <= 9'b11110101;
				8'b101101: c <= 9'b10111001;
				8'b1010011: c <= 9'b11001110;
				8'b1100001: c <= 9'b111001;
				8'b110101: c <= 9'b1111010;
				8'b1000100: c <= 9'b101110001;
				8'b1010001: c <= 9'b111111111;
				8'b1010100: c <= 9'b110111000;
				8'b1100110: c <= 9'b110010100;
				8'b101010: c <= 9'b100110000;
				8'b1011110: c <= 9'b11000100;
				8'b1100111: c <= 9'b1100011;
				8'b1011010: c <= 9'b10011010;
				8'b1000010: c <= 9'b111101;
				8'b111101: c <= 9'b101111111;
				8'b110000: c <= 9'b111111011;
				8'b111110: c <= 9'b101100010;
				8'b1100010: c <= 9'b101100;
				8'b1110000: c <= 9'b11100000;
				8'b1101001: c <= 9'b101001;
				8'b1110011: c <= 9'b11110;
				8'b1001100: c <= 9'b100;
				8'b100001: c <= 9'b11011000;
				8'b1000110: c <= 9'b100101110;
				8'b1110010: c <= 9'b110001111;
				8'b1010000: c <= 9'b1110100;
				8'b1111010: c <= 9'b100110010;
				8'b1010101: c <= 9'b100011001;
				8'b111011: c <= 9'b1011000;
				8'b1001101: c <= 9'b110111000;
				8'b111111: c <= 9'b1000111;
				8'b1101110: c <= 9'b11000110;
				8'b1111011: c <= 9'b11001;
				8'b1001011: c <= 9'b100011000;
				8'b1101111: c <= 9'b101101110;
				8'b1101000: c <= 9'b100010001;
				8'b101100: c <= 9'b101100111;
				8'b100100: c <= 9'b11011;
				8'b1111000: c <= 9'b10011100;
				8'b1000101: c <= 9'b10001010;
				8'b1011001: c <= 9'b101010000;
				8'b110100: c <= 9'b11011001;
				8'b1111001: c <= 9'b10011101;
				8'b1110001: c <= 9'b111001;
				8'b1001111: c <= 9'b101;
				8'b1100101: c <= 9'b100000010;
				8'b1111110: c <= 9'b111001101;
				8'b1111100: c <= 9'b10101;
				8'b1010110: c <= 9'b110111111;
				8'b110010: c <= 9'b11000000;
				8'b1101101: c <= 9'b111101110;
				8'b100011: c <= 9'b100001;
				8'b1110101: c <= 9'b11100000;
				8'b1111101: c <= 9'b110001000;
				8'b101001: c <= 9'b11101111;
				8'b1010010: c <= 9'b10010;
				8'b1011000: c <= 9'b100101111;
				8'b101110: c <= 9'b10111101;
				8'b1000001: c <= 9'b100110010;
				default: c <= 9'b0;
			endcase
			9'b10111100 : case(di)
				8'b1000011: c <= 9'b111000111;
				8'b101000: c <= 9'b110000101;
				8'b111010: c <= 9'b111011010;
				8'b110110: c <= 9'b101010;
				8'b1100100: c <= 9'b111010111;
				8'b1000000: c <= 9'b11001001;
				8'b1110110: c <= 9'b110001001;
				8'b100101: c <= 9'b11;
				8'b101111: c <= 9'b10111010;
				8'b100110: c <= 9'b110100110;
				8'b1100011: c <= 9'b1111111;
				8'b1001000: c <= 9'b110101101;
				8'b111000: c <= 9'b10011101;
				8'b110001: c <= 9'b110000010;
				8'b1010111: c <= 9'b111011100;
				8'b1001110: c <= 9'b101000101;
				8'b1101010: c <= 9'b100100011;
				8'b1001001: c <= 9'b100000100;
				8'b1100000: c <= 9'b10101010;
				8'b110111: c <= 9'b11111010;
				8'b1011101: c <= 9'b111001011;
				8'b1011011: c <= 9'b10100010;
				8'b111001: c <= 9'b111110001;
				8'b1001010: c <= 9'b110010010;
				8'b110011: c <= 9'b110100000;
				8'b1101100: c <= 9'b10011111;
				8'b1110111: c <= 9'b111101110;
				8'b101011: c <= 9'b1100000;
				8'b1101011: c <= 9'b110111100;
				8'b111100: c <= 9'b1111011;
				8'b1000111: c <= 9'b110011011;
				8'b1011111: c <= 9'b100101111;
				8'b1110100: c <= 9'b110100;
				8'b101101: c <= 9'b100011011;
				8'b1010011: c <= 9'b100010000;
				8'b1100001: c <= 9'b10101000;
				8'b110101: c <= 9'b110011110;
				8'b1000100: c <= 9'b111100101;
				8'b1010001: c <= 9'b10000011;
				8'b1010100: c <= 9'b11010101;
				8'b1100110: c <= 9'b100110111;
				8'b101010: c <= 9'b111000101;
				8'b1011110: c <= 9'b11111100;
				8'b1100111: c <= 9'b11110001;
				8'b1011010: c <= 9'b101001;
				8'b1000010: c <= 9'b111110011;
				8'b111101: c <= 9'b10100010;
				8'b110000: c <= 9'b1000001;
				8'b111110: c <= 9'b110010011;
				8'b1100010: c <= 9'b110111011;
				8'b1110000: c <= 9'b100111000;
				8'b1101001: c <= 9'b101101000;
				8'b1110011: c <= 9'b110100;
				8'b1001100: c <= 9'b100110011;
				8'b100001: c <= 9'b100111011;
				8'b1000110: c <= 9'b110110010;
				8'b1110010: c <= 9'b10101111;
				8'b1010000: c <= 9'b111111011;
				8'b1111010: c <= 9'b111100001;
				8'b1010101: c <= 9'b110011000;
				8'b111011: c <= 9'b110100101;
				8'b1001101: c <= 9'b100001101;
				8'b111111: c <= 9'b111000100;
				8'b1101110: c <= 9'b11110001;
				8'b1111011: c <= 9'b11011011;
				8'b1001011: c <= 9'b111011010;
				8'b1101111: c <= 9'b101001110;
				8'b1101000: c <= 9'b11100;
				8'b101100: c <= 9'b10010111;
				8'b100100: c <= 9'b1111010;
				8'b1111000: c <= 9'b101101001;
				8'b1000101: c <= 9'b1110100;
				8'b1011001: c <= 9'b1001000;
				8'b110100: c <= 9'b111111000;
				8'b1111001: c <= 9'b110010;
				8'b1110001: c <= 9'b10100010;
				8'b1001111: c <= 9'b1;
				8'b1100101: c <= 9'b110101010;
				8'b1111110: c <= 9'b1100;
				8'b1111100: c <= 9'b10110011;
				8'b1010110: c <= 9'b101001111;
				8'b110010: c <= 9'b1001001;
				8'b1101101: c <= 9'b11111100;
				8'b100011: c <= 9'b11100111;
				8'b1110101: c <= 9'b11100011;
				8'b1111101: c <= 9'b110011111;
				8'b101001: c <= 9'b101111010;
				8'b1010010: c <= 9'b1010000;
				8'b1011000: c <= 9'b100001111;
				8'b101110: c <= 9'b100101010;
				8'b1000001: c <= 9'b110000110;
				default: c <= 9'b0;
			endcase
			9'b10101011 : case(di)
				8'b1000011: c <= 9'b111101000;
				8'b101000: c <= 9'b101011;
				8'b111010: c <= 9'b110100111;
				8'b110110: c <= 9'b110100001;
				8'b1100100: c <= 9'b10010110;
				8'b1000000: c <= 9'b100101;
				8'b1110110: c <= 9'b101001000;
				8'b100101: c <= 9'b110000111;
				8'b101111: c <= 9'b100101110;
				8'b100110: c <= 9'b10100101;
				8'b1100011: c <= 9'b101001010;
				8'b1001000: c <= 9'b111111110;
				8'b111000: c <= 9'b100101011;
				8'b110001: c <= 9'b10000011;
				8'b1010111: c <= 9'b100100010;
				8'b1001110: c <= 9'b10100010;
				8'b1101010: c <= 9'b11011011;
				8'b1001001: c <= 9'b111100011;
				8'b1100000: c <= 9'b1001001;
				8'b110111: c <= 9'b100001001;
				8'b1011101: c <= 9'b10100;
				8'b1011011: c <= 9'b101010110;
				8'b111001: c <= 9'b100011;
				8'b1001010: c <= 9'b110111001;
				8'b110011: c <= 9'b10;
				8'b1101100: c <= 9'b110001010;
				8'b1110111: c <= 9'b100;
				8'b101011: c <= 9'b110100100;
				8'b1101011: c <= 9'b111101110;
				8'b111100: c <= 9'b101000;
				8'b1000111: c <= 9'b110111011;
				8'b1011111: c <= 9'b1110101;
				8'b1110100: c <= 9'b101000011;
				8'b101101: c <= 9'b11011010;
				8'b1010011: c <= 9'b100110100;
				8'b1100001: c <= 9'b110000;
				8'b110101: c <= 9'b110100001;
				8'b1000100: c <= 9'b1001101;
				8'b1010001: c <= 9'b100101111;
				8'b1010100: c <= 9'b110110011;
				8'b1100110: c <= 9'b110011001;
				8'b101010: c <= 9'b110000110;
				8'b1011110: c <= 9'b101111001;
				8'b1100111: c <= 9'b101000111;
				8'b1011010: c <= 9'b1000010;
				8'b1000010: c <= 9'b10111100;
				8'b111101: c <= 9'b10100111;
				8'b110000: c <= 9'b110100101;
				8'b111110: c <= 9'b101001100;
				8'b1100010: c <= 9'b10000011;
				8'b1110000: c <= 9'b110000011;
				8'b1101001: c <= 9'b11100100;
				8'b1110011: c <= 9'b11000011;
				8'b1001100: c <= 9'b100101001;
				8'b100001: c <= 9'b110111110;
				8'b1000110: c <= 9'b1110010;
				8'b1110010: c <= 9'b10010001;
				8'b1010000: c <= 9'b111001111;
				8'b1111010: c <= 9'b1011001;
				8'b1010101: c <= 9'b100000101;
				8'b111011: c <= 9'b1111011;
				8'b1001101: c <= 9'b100111000;
				8'b111111: c <= 9'b101010110;
				8'b1101110: c <= 9'b101010001;
				8'b1111011: c <= 9'b11110101;
				8'b1001011: c <= 9'b101000101;
				8'b1101111: c <= 9'b110001;
				8'b1101000: c <= 9'b1010010;
				8'b101100: c <= 9'b1000;
				8'b100100: c <= 9'b110100100;
				8'b1111000: c <= 9'b1011;
				8'b1000101: c <= 9'b1100011;
				8'b1011001: c <= 9'b1000101;
				8'b110100: c <= 9'b100101110;
				8'b1111001: c <= 9'b100010111;
				8'b1110001: c <= 9'b110000011;
				8'b1001111: c <= 9'b111100000;
				8'b1100101: c <= 9'b11001110;
				8'b1111110: c <= 9'b10101000;
				8'b1111100: c <= 9'b11101101;
				8'b1010110: c <= 9'b11001;
				8'b110010: c <= 9'b110010;
				8'b1101101: c <= 9'b110010100;
				8'b100011: c <= 9'b1000110;
				8'b1110101: c <= 9'b110110010;
				8'b1111101: c <= 9'b111101110;
				8'b101001: c <= 9'b10110101;
				8'b1010010: c <= 9'b110000101;
				8'b1011000: c <= 9'b110111001;
				8'b101110: c <= 9'b100010;
				8'b1000001: c <= 9'b110011100;
				default: c <= 9'b0;
			endcase
			9'b11110001 : case(di)
				8'b1000011: c <= 9'b111001001;
				8'b101000: c <= 9'b110101110;
				8'b111010: c <= 9'b101000110;
				8'b110110: c <= 9'b10110001;
				8'b1100100: c <= 9'b111001101;
				8'b1000000: c <= 9'b100101101;
				8'b1110110: c <= 9'b10101011;
				8'b100101: c <= 9'b1110111;
				8'b101111: c <= 9'b111001110;
				8'b100110: c <= 9'b110010101;
				8'b1100011: c <= 9'b1110000;
				8'b1001000: c <= 9'b110110110;
				8'b111000: c <= 9'b100100010;
				8'b110001: c <= 9'b100010111;
				8'b1010111: c <= 9'b100000000;
				8'b1001110: c <= 9'b100101101;
				8'b1101010: c <= 9'b101011000;
				8'b1001001: c <= 9'b10010000;
				8'b1100000: c <= 9'b111100100;
				8'b110111: c <= 9'b111001;
				8'b1011101: c <= 9'b1100110;
				8'b1011011: c <= 9'b101111010;
				8'b111001: c <= 9'b100001110;
				8'b1001010: c <= 9'b101000110;
				8'b110011: c <= 9'b11110011;
				8'b1101100: c <= 9'b110010110;
				8'b1110111: c <= 9'b101010100;
				8'b101011: c <= 9'b110001000;
				8'b1101011: c <= 9'b110010110;
				8'b111100: c <= 9'b101110001;
				8'b1000111: c <= 9'b11010001;
				8'b1011111: c <= 9'b111101000;
				8'b1110100: c <= 9'b101101010;
				8'b101101: c <= 9'b10100010;
				8'b1010011: c <= 9'b11000100;
				8'b1100001: c <= 9'b10101001;
				8'b110101: c <= 9'b100001100;
				8'b1000100: c <= 9'b110100000;
				8'b1010001: c <= 9'b1010010;
				8'b1010100: c <= 9'b111101111;
				8'b1100110: c <= 9'b100111;
				8'b101010: c <= 9'b101001011;
				8'b1011110: c <= 9'b11101101;
				8'b1100111: c <= 9'b110010;
				8'b1011010: c <= 9'b111001010;
				8'b1000010: c <= 9'b1110100;
				8'b111101: c <= 9'b100001100;
				8'b110000: c <= 9'b100111010;
				8'b111110: c <= 9'b110100111;
				8'b1100010: c <= 9'b101101110;
				8'b1110000: c <= 9'b100011011;
				8'b1101001: c <= 9'b10110011;
				8'b1110011: c <= 9'b1000011;
				8'b1001100: c <= 9'b11100101;
				8'b100001: c <= 9'b110000001;
				8'b1000110: c <= 9'b100010111;
				8'b1110010: c <= 9'b110110000;
				8'b1010000: c <= 9'b100011000;
				8'b1111010: c <= 9'b1111;
				8'b1010101: c <= 9'b101101111;
				8'b111011: c <= 9'b11100010;
				8'b1001101: c <= 9'b1000100;
				8'b111111: c <= 9'b110111011;
				8'b1101110: c <= 9'b101001011;
				8'b1111011: c <= 9'b1011100;
				8'b1001011: c <= 9'b10100000;
				8'b1101111: c <= 9'b1000;
				8'b1101000: c <= 9'b100011100;
				8'b101100: c <= 9'b110110;
				8'b100100: c <= 9'b10101001;
				8'b1111000: c <= 9'b110101101;
				8'b1000101: c <= 9'b1010001;
				8'b1011001: c <= 9'b110101;
				8'b110100: c <= 9'b101000011;
				8'b1111001: c <= 9'b100101000;
				8'b1110001: c <= 9'b110111100;
				8'b1001111: c <= 9'b11110011;
				8'b1100101: c <= 9'b111111001;
				8'b1111110: c <= 9'b111000000;
				8'b1111100: c <= 9'b111101000;
				8'b1010110: c <= 9'b10001010;
				8'b110010: c <= 9'b11111011;
				8'b1101101: c <= 9'b100001;
				8'b100011: c <= 9'b110110;
				8'b1110101: c <= 9'b101100001;
				8'b1111101: c <= 9'b100111100;
				8'b101001: c <= 9'b100000010;
				8'b1010010: c <= 9'b101110010;
				8'b1011000: c <= 9'b10011000;
				8'b101110: c <= 9'b101101;
				8'b1000001: c <= 9'b1100111;
				default: c <= 9'b0;
			endcase
			9'b11000 : case(di)
				8'b1000011: c <= 9'b11110100;
				8'b101000: c <= 9'b1111001;
				8'b111010: c <= 9'b11111011;
				8'b110110: c <= 9'b10000001;
				8'b1100100: c <= 9'b10010011;
				8'b1000000: c <= 9'b100101111;
				8'b1110110: c <= 9'b101001001;
				8'b100101: c <= 9'b100101111;
				8'b101111: c <= 9'b100011100;
				8'b100110: c <= 9'b110010011;
				8'b1100011: c <= 9'b101101010;
				8'b1001000: c <= 9'b110010010;
				8'b111000: c <= 9'b100101001;
				8'b110001: c <= 9'b100100001;
				8'b1010111: c <= 9'b101011110;
				8'b1001110: c <= 9'b1100100;
				8'b1101010: c <= 9'b1101001;
				8'b1001001: c <= 9'b100011010;
				8'b1100000: c <= 9'b101010100;
				8'b110111: c <= 9'b110111011;
				8'b1011101: c <= 9'b1001110;
				8'b1011011: c <= 9'b10010111;
				8'b111001: c <= 9'b11010011;
				8'b1001010: c <= 9'b110100100;
				8'b110011: c <= 9'b101000011;
				8'b1101100: c <= 9'b110001000;
				8'b1110111: c <= 9'b101001;
				8'b101011: c <= 9'b100001010;
				8'b1101011: c <= 9'b11000;
				8'b111100: c <= 9'b11001101;
				8'b1000111: c <= 9'b100111000;
				8'b1011111: c <= 9'b10010111;
				8'b1110100: c <= 9'b110001;
				8'b101101: c <= 9'b111010010;
				8'b1010011: c <= 9'b11011100;
				8'b1100001: c <= 9'b111100000;
				8'b110101: c <= 9'b101011011;
				8'b1000100: c <= 9'b100011100;
				8'b1010001: c <= 9'b10100111;
				8'b1010100: c <= 9'b101010000;
				8'b1100110: c <= 9'b101100010;
				8'b101010: c <= 9'b110011001;
				8'b1011110: c <= 9'b1010111;
				8'b1100111: c <= 9'b111001;
				8'b1011010: c <= 9'b101001;
				8'b1000010: c <= 9'b111000010;
				8'b111101: c <= 9'b110011010;
				8'b110000: c <= 9'b1100111;
				8'b111110: c <= 9'b110100;
				8'b1100010: c <= 9'b111100;
				8'b1110000: c <= 9'b110101;
				8'b1101001: c <= 9'b11111010;
				8'b1110011: c <= 9'b110101101;
				8'b1001100: c <= 9'b10111111;
				8'b100001: c <= 9'b111010010;
				8'b1000110: c <= 9'b101100001;
				8'b1110010: c <= 9'b10110001;
				8'b1010000: c <= 9'b11101101;
				8'b1111010: c <= 9'b101110000;
				8'b1010101: c <= 9'b110000;
				8'b111011: c <= 9'b101100101;
				8'b1001101: c <= 9'b100011000;
				8'b111111: c <= 9'b1111110;
				8'b1101110: c <= 9'b100;
				8'b1111011: c <= 9'b1010101;
				8'b1001011: c <= 9'b1111011;
				8'b1101111: c <= 9'b101110010;
				8'b1101000: c <= 9'b100101110;
				8'b101100: c <= 9'b100001101;
				8'b100100: c <= 9'b1111101;
				8'b1111000: c <= 9'b100000001;
				8'b1000101: c <= 9'b100;
				8'b1011001: c <= 9'b110001110;
				8'b110100: c <= 9'b10010110;
				8'b1111001: c <= 9'b111001111;
				8'b1110001: c <= 9'b110001010;
				8'b1001111: c <= 9'b101010;
				8'b1100101: c <= 9'b101011110;
				8'b1111110: c <= 9'b10111000;
				8'b1111100: c <= 9'b10001110;
				8'b1010110: c <= 9'b110101010;
				8'b110010: c <= 9'b11110010;
				8'b1101101: c <= 9'b11010001;
				8'b100011: c <= 9'b101001110;
				8'b1110101: c <= 9'b1000110;
				8'b1111101: c <= 9'b100010111;
				8'b101001: c <= 9'b11100101;
				8'b1010010: c <= 9'b110111011;
				8'b1011000: c <= 9'b101000;
				8'b101110: c <= 9'b1001110;
				8'b1000001: c <= 9'b1001111;
				default: c <= 9'b0;
			endcase
			9'b11000010 : case(di)
				8'b1000011: c <= 9'b111010010;
				8'b101000: c <= 9'b110100001;
				8'b111010: c <= 9'b110000;
				8'b110110: c <= 9'b11;
				8'b1100100: c <= 9'b110111100;
				8'b1000000: c <= 9'b101100110;
				8'b1110110: c <= 9'b111111001;
				8'b100101: c <= 9'b1001000;
				8'b101111: c <= 9'b110101011;
				8'b100110: c <= 9'b1100101;
				8'b1100011: c <= 9'b1101100;
				8'b1001000: c <= 9'b111100001;
				8'b111000: c <= 9'b110111011;
				8'b110001: c <= 9'b10101000;
				8'b1010111: c <= 9'b111101110;
				8'b1001110: c <= 9'b111111;
				8'b1101010: c <= 9'b10110100;
				8'b1001001: c <= 9'b110010101;
				8'b1100000: c <= 9'b1100010;
				8'b110111: c <= 9'b100100;
				8'b1011101: c <= 9'b10100101;
				8'b1011011: c <= 9'b110000111;
				8'b111001: c <= 9'b101010;
				8'b1001010: c <= 9'b110110010;
				8'b110011: c <= 9'b111100011;
				8'b1101100: c <= 9'b110100011;
				8'b1110111: c <= 9'b11101111;
				8'b101011: c <= 9'b101000;
				8'b1101011: c <= 9'b111001100;
				8'b111100: c <= 9'b11000110;
				8'b1000111: c <= 9'b1000101;
				8'b1011111: c <= 9'b101000011;
				8'b1110100: c <= 9'b110001101;
				8'b101101: c <= 9'b100110111;
				8'b1010011: c <= 9'b1011;
				8'b1100001: c <= 9'b1110010;
				8'b110101: c <= 9'b110111011;
				8'b1000100: c <= 9'b101110001;
				8'b1010001: c <= 9'b1001110;
				8'b1010100: c <= 9'b101011101;
				8'b1100110: c <= 9'b100101011;
				8'b101010: c <= 9'b100100111;
				8'b1011110: c <= 9'b1010010;
				8'b1100111: c <= 9'b100011010;
				8'b1011010: c <= 9'b111010111;
				8'b1000010: c <= 9'b101101111;
				8'b111101: c <= 9'b111101111;
				8'b110000: c <= 9'b1001101;
				8'b111110: c <= 9'b10000011;
				8'b1100010: c <= 9'b11010;
				8'b1110000: c <= 9'b101000001;
				8'b1101001: c <= 9'b111000;
				8'b1110011: c <= 9'b111110000;
				8'b1001100: c <= 9'b101010010;
				8'b100001: c <= 9'b110101110;
				8'b1000110: c <= 9'b111100100;
				8'b1110010: c <= 9'b11001100;
				8'b1010000: c <= 9'b100100011;
				8'b1111010: c <= 9'b10010;
				8'b1010101: c <= 9'b110100110;
				8'b111011: c <= 9'b1110111;
				8'b1001101: c <= 9'b101111001;
				8'b111111: c <= 9'b110001111;
				8'b1101110: c <= 9'b110011010;
				8'b1111011: c <= 9'b11000000;
				8'b1001011: c <= 9'b1010011;
				8'b1101111: c <= 9'b100100000;
				8'b1101000: c <= 9'b101100001;
				8'b101100: c <= 9'b10111111;
				8'b100100: c <= 9'b110010;
				8'b1111000: c <= 9'b100011001;
				8'b1000101: c <= 9'b111011;
				8'b1011001: c <= 9'b111111011;
				8'b110100: c <= 9'b111001010;
				8'b1111001: c <= 9'b111101100;
				8'b1110001: c <= 9'b100000111;
				8'b1001111: c <= 9'b10010100;
				8'b1100101: c <= 9'b111111011;
				8'b1111110: c <= 9'b100111111;
				8'b1111100: c <= 9'b111011001;
				8'b1010110: c <= 9'b110100010;
				8'b110010: c <= 9'b10001001;
				8'b1101101: c <= 9'b110011110;
				8'b100011: c <= 9'b110000011;
				8'b1110101: c <= 9'b11100101;
				8'b1111101: c <= 9'b111011101;
				8'b101001: c <= 9'b1010110;
				8'b1010010: c <= 9'b1011011;
				8'b1011000: c <= 9'b1110011;
				8'b101110: c <= 9'b1000011;
				8'b1000001: c <= 9'b11100100;
				default: c <= 9'b0;
			endcase
			9'b100000101 : case(di)
				8'b1000011: c <= 9'b10100111;
				8'b101000: c <= 9'b101000101;
				8'b111010: c <= 9'b100100011;
				8'b110110: c <= 9'b100000000;
				8'b1100100: c <= 9'b100110011;
				8'b1000000: c <= 9'b100100001;
				8'b1110110: c <= 9'b11011001;
				8'b100101: c <= 9'b110010010;
				8'b101111: c <= 9'b1000000;
				8'b100110: c <= 9'b101010110;
				8'b1100011: c <= 9'b110;
				8'b1001000: c <= 9'b1000;
				8'b111000: c <= 9'b111110110;
				8'b110001: c <= 9'b11000011;
				8'b1010111: c <= 9'b111100101;
				8'b1001110: c <= 9'b10010100;
				8'b1101010: c <= 9'b10101101;
				8'b1001001: c <= 9'b1010111;
				8'b1100000: c <= 9'b101110;
				8'b110111: c <= 9'b10101;
				8'b1011101: c <= 9'b101100000;
				8'b1011011: c <= 9'b111101000;
				8'b111001: c <= 9'b11111010;
				8'b1001010: c <= 9'b11111010;
				8'b110011: c <= 9'b100000101;
				8'b1101100: c <= 9'b1101000;
				8'b1110111: c <= 9'b110001011;
				8'b101011: c <= 9'b1000;
				8'b1101011: c <= 9'b11101101;
				8'b111100: c <= 9'b11111010;
				8'b1000111: c <= 9'b11011001;
				8'b1011111: c <= 9'b110101110;
				8'b1110100: c <= 9'b101000011;
				8'b101101: c <= 9'b101001110;
				8'b1010011: c <= 9'b111000010;
				8'b1100001: c <= 9'b100001100;
				8'b110101: c <= 9'b10010011;
				8'b1000100: c <= 9'b110011;
				8'b1010001: c <= 9'b1110011;
				8'b1010100: c <= 9'b1110;
				8'b1100110: c <= 9'b101110001;
				8'b101010: c <= 9'b11011110;
				8'b1011110: c <= 9'b11100111;
				8'b1100111: c <= 9'b101010011;
				8'b1011010: c <= 9'b101001;
				8'b1000010: c <= 9'b100110;
				8'b111101: c <= 9'b110000001;
				8'b110000: c <= 9'b11010001;
				8'b111110: c <= 9'b100000000;
				8'b1100010: c <= 9'b101010000;
				8'b1110000: c <= 9'b11000001;
				8'b1101001: c <= 9'b101001110;
				8'b1110011: c <= 9'b101111010;
				8'b1001100: c <= 9'b1101110;
				8'b100001: c <= 9'b11010001;
				8'b1000110: c <= 9'b101101011;
				8'b1110010: c <= 9'b100100010;
				8'b1010000: c <= 9'b101011001;
				8'b1111010: c <= 9'b100001100;
				8'b1010101: c <= 9'b11010111;
				8'b111011: c <= 9'b1001000;
				8'b1001101: c <= 9'b110011100;
				8'b111111: c <= 9'b11011001;
				8'b1101110: c <= 9'b101011000;
				8'b1111011: c <= 9'b1001000;
				8'b1001011: c <= 9'b100011;
				8'b1101111: c <= 9'b11011100;
				8'b1101000: c <= 9'b101110001;
				8'b101100: c <= 9'b100101010;
				8'b100100: c <= 9'b100111011;
				8'b1111000: c <= 9'b11111100;
				8'b1000101: c <= 9'b100001001;
				8'b1011001: c <= 9'b101100110;
				8'b110100: c <= 9'b100011111;
				8'b1111001: c <= 9'b101010;
				8'b1110001: c <= 9'b101001111;
				8'b1001111: c <= 9'b111000011;
				8'b1100101: c <= 9'b100100011;
				8'b1111110: c <= 9'b100110010;
				8'b1111100: c <= 9'b100001010;
				8'b1010110: c <= 9'b111101111;
				8'b110010: c <= 9'b111101111;
				8'b1101101: c <= 9'b100100;
				8'b100011: c <= 9'b100000111;
				8'b1110101: c <= 9'b110110100;
				8'b1111101: c <= 9'b100010100;
				8'b101001: c <= 9'b1111111;
				8'b1010010: c <= 9'b1110001;
				8'b1011000: c <= 9'b10011100;
				8'b101110: c <= 9'b11010111;
				8'b1000001: c <= 9'b1010110;
				default: c <= 9'b0;
			endcase
			9'b100111100 : case(di)
				8'b1000011: c <= 9'b110001001;
				8'b101000: c <= 9'b11011000;
				8'b111010: c <= 9'b110011010;
				8'b110110: c <= 9'b1110010;
				8'b1100100: c <= 9'b10001100;
				8'b1000000: c <= 9'b100000101;
				8'b1110110: c <= 9'b101000010;
				8'b100101: c <= 9'b100001001;
				8'b101111: c <= 9'b10101010;
				8'b100110: c <= 9'b110011110;
				8'b1100011: c <= 9'b1111000;
				8'b1001000: c <= 9'b100011;
				8'b111000: c <= 9'b111000101;
				8'b110001: c <= 9'b110001110;
				8'b1010111: c <= 9'b100100000;
				8'b1001110: c <= 9'b101000111;
				8'b1101010: c <= 9'b101010110;
				8'b1001001: c <= 9'b110111111;
				8'b1100000: c <= 9'b101010010;
				8'b110111: c <= 9'b1010111;
				8'b1011101: c <= 9'b10101;
				8'b1011011: c <= 9'b110100110;
				8'b111001: c <= 9'b11010100;
				8'b1001010: c <= 9'b1110101;
				8'b110011: c <= 9'b100000101;
				8'b1101100: c <= 9'b11101100;
				8'b1110111: c <= 9'b10001100;
				8'b101011: c <= 9'b101110101;
				8'b1101011: c <= 9'b1110011;
				8'b111100: c <= 9'b111100;
				8'b1000111: c <= 9'b10101010;
				8'b1011111: c <= 9'b101001010;
				8'b1110100: c <= 9'b100110100;
				8'b101101: c <= 9'b100100;
				8'b1010011: c <= 9'b101111110;
				8'b1100001: c <= 9'b100111000;
				8'b110101: c <= 9'b101110010;
				8'b1000100: c <= 9'b1010010;
				8'b1010001: c <= 9'b1000011;
				8'b1010100: c <= 9'b11100111;
				8'b1100110: c <= 9'b101011;
				8'b101010: c <= 9'b11111010;
				8'b1011110: c <= 9'b101110000;
				8'b1100111: c <= 9'b111000111;
				8'b1011010: c <= 9'b11001000;
				8'b1000010: c <= 9'b10100111;
				8'b111101: c <= 9'b10100100;
				8'b110000: c <= 9'b111101000;
				8'b111110: c <= 9'b111100111;
				8'b1100010: c <= 9'b111111010;
				8'b1110000: c <= 9'b1111110;
				8'b1101001: c <= 9'b100011111;
				8'b1110011: c <= 9'b110010;
				8'b1001100: c <= 9'b101110000;
				8'b100001: c <= 9'b101100;
				8'b1000110: c <= 9'b11000;
				8'b1110010: c <= 9'b10110100;
				8'b1010000: c <= 9'b111111111;
				8'b1111010: c <= 9'b110000010;
				8'b1010101: c <= 9'b10011001;
				8'b111011: c <= 9'b111011010;
				8'b1001101: c <= 9'b10101;
				8'b111111: c <= 9'b10;
				8'b1101110: c <= 9'b111110000;
				8'b1111011: c <= 9'b100001;
				8'b1001011: c <= 9'b11000111;
				8'b1101111: c <= 9'b1110000;
				8'b1101000: c <= 9'b1101000;
				8'b101100: c <= 9'b100011111;
				8'b100100: c <= 9'b110111000;
				8'b1111000: c <= 9'b110100110;
				8'b1000101: c <= 9'b111110001;
				8'b1011001: c <= 9'b110000110;
				8'b110100: c <= 9'b10100011;
				8'b1111001: c <= 9'b10111110;
				8'b1110001: c <= 9'b111000000;
				8'b1001111: c <= 9'b11011100;
				8'b1100101: c <= 9'b101011001;
				8'b1111110: c <= 9'b101111000;
				8'b1111100: c <= 9'b100100;
				8'b1010110: c <= 9'b1011111;
				8'b110010: c <= 9'b10110111;
				8'b1101101: c <= 9'b11111000;
				8'b100011: c <= 9'b111011101;
				8'b1110101: c <= 9'b101001111;
				8'b1111101: c <= 9'b111001110;
				8'b101001: c <= 9'b100111110;
				8'b1010010: c <= 9'b10111000;
				8'b1011000: c <= 9'b10010001;
				8'b101110: c <= 9'b100010000;
				8'b1000001: c <= 9'b11000110;
				default: c <= 9'b0;
			endcase
			9'b111110001 : case(di)
				8'b1000011: c <= 9'b100011000;
				8'b101000: c <= 9'b1110101;
				8'b111010: c <= 9'b1111011;
				8'b110110: c <= 9'b1110010;
				8'b1100100: c <= 9'b101111001;
				8'b1000000: c <= 9'b11011101;
				8'b1110110: c <= 9'b111111110;
				8'b100101: c <= 9'b111111011;
				8'b101111: c <= 9'b100100111;
				8'b100110: c <= 9'b10100110;
				8'b1100011: c <= 9'b11000;
				8'b1001000: c <= 9'b1111011;
				8'b111000: c <= 9'b1;
				8'b110001: c <= 9'b100010111;
				8'b1010111: c <= 9'b100111011;
				8'b1001110: c <= 9'b100110;
				8'b1101010: c <= 9'b100110101;
				8'b1001001: c <= 9'b11000000;
				8'b1100000: c <= 9'b110110100;
				8'b110111: c <= 9'b101110111;
				8'b1011101: c <= 9'b1110;
				8'b1011011: c <= 9'b111000000;
				8'b111001: c <= 9'b101011000;
				8'b1001010: c <= 9'b111001;
				8'b110011: c <= 9'b100000110;
				8'b1101100: c <= 9'b10011;
				8'b1110111: c <= 9'b10101101;
				8'b101011: c <= 9'b10001010;
				8'b1101011: c <= 9'b1100000;
				8'b111100: c <= 9'b100010001;
				8'b1000111: c <= 9'b11110100;
				8'b1011111: c <= 9'b1001001;
				8'b1110100: c <= 9'b100000111;
				8'b101101: c <= 9'b11111010;
				8'b1010011: c <= 9'b110100101;
				8'b1100001: c <= 9'b11101011;
				8'b110101: c <= 9'b1101101;
				8'b1000100: c <= 9'b111100101;
				8'b1010001: c <= 9'b101110011;
				8'b1010100: c <= 9'b110101111;
				8'b1100110: c <= 9'b100010;
				8'b101010: c <= 9'b101100001;
				8'b1011110: c <= 9'b110111110;
				8'b1100111: c <= 9'b1110;
				8'b1011010: c <= 9'b101100;
				8'b1000010: c <= 9'b111001011;
				8'b111101: c <= 9'b101100100;
				8'b110000: c <= 9'b110000001;
				8'b111110: c <= 9'b111001111;
				8'b1100010: c <= 9'b100110100;
				8'b1110000: c <= 9'b10111011;
				8'b1101001: c <= 9'b111111111;
				8'b1110011: c <= 9'b111000111;
				8'b1001100: c <= 9'b100000001;
				8'b100001: c <= 9'b101110000;
				8'b1000110: c <= 9'b100011101;
				8'b1110010: c <= 9'b100010101;
				8'b1010000: c <= 9'b10001110;
				8'b1111010: c <= 9'b110101011;
				8'b1010101: c <= 9'b10110110;
				8'b111011: c <= 9'b101101110;
				8'b1001101: c <= 9'b11111001;
				8'b111111: c <= 9'b1110;
				8'b1101110: c <= 9'b101110001;
				8'b1111011: c <= 9'b111010111;
				8'b1001011: c <= 9'b1001000;
				8'b1101111: c <= 9'b100101010;
				8'b1101000: c <= 9'b11010001;
				8'b101100: c <= 9'b10110111;
				8'b100100: c <= 9'b101011010;
				8'b1111000: c <= 9'b100010000;
				8'b1000101: c <= 9'b100111111;
				8'b1011001: c <= 9'b111010110;
				8'b110100: c <= 9'b1001;
				8'b1111001: c <= 9'b100001011;
				8'b1110001: c <= 9'b11111001;
				8'b1001111: c <= 9'b100110010;
				8'b1100101: c <= 9'b11100101;
				8'b1111110: c <= 9'b11101100;
				8'b1111100: c <= 9'b110111111;
				8'b1010110: c <= 9'b11000;
				8'b110010: c <= 9'b101101110;
				8'b1101101: c <= 9'b1000;
				8'b100011: c <= 9'b10;
				8'b1110101: c <= 9'b110010111;
				8'b1111101: c <= 9'b10000110;
				8'b101001: c <= 9'b111110110;
				8'b1010010: c <= 9'b111010110;
				8'b1011000: c <= 9'b101101111;
				8'b101110: c <= 9'b1101101;
				8'b1000001: c <= 9'b10101110;
				default: c <= 9'b0;
			endcase
			9'b100100 : case(di)
				8'b1000011: c <= 9'b111010110;
				8'b101000: c <= 9'b10010111;
				8'b111010: c <= 9'b111100111;
				8'b110110: c <= 9'b111010111;
				8'b1100100: c <= 9'b101110100;
				8'b1000000: c <= 9'b1011000;
				8'b1110110: c <= 9'b101011110;
				8'b100101: c <= 9'b11110010;
				8'b101111: c <= 9'b110011101;
				8'b100110: c <= 9'b110001110;
				8'b1100011: c <= 9'b101101001;
				8'b1001000: c <= 9'b1001011;
				8'b111000: c <= 9'b111011010;
				8'b110001: c <= 9'b110101011;
				8'b1010111: c <= 9'b1011001;
				8'b1001110: c <= 9'b10011111;
				8'b1101010: c <= 9'b11001000;
				8'b1001001: c <= 9'b110100011;
				8'b1100000: c <= 9'b10110011;
				8'b110111: c <= 9'b100001;
				8'b1011101: c <= 9'b101011111;
				8'b1011011: c <= 9'b11000001;
				8'b111001: c <= 9'b100010010;
				8'b1001010: c <= 9'b10111100;
				8'b110011: c <= 9'b110101011;
				8'b1101100: c <= 9'b100101110;
				8'b1110111: c <= 9'b11010010;
				8'b101011: c <= 9'b100000001;
				8'b1101011: c <= 9'b1010001;
				8'b111100: c <= 9'b100001111;
				8'b1000111: c <= 9'b110001110;
				8'b1011111: c <= 9'b1010000;
				8'b1110100: c <= 9'b11000111;
				8'b101101: c <= 9'b11100000;
				8'b1010011: c <= 9'b11100001;
				8'b1100001: c <= 9'b101110;
				8'b110101: c <= 9'b110111110;
				8'b1000100: c <= 9'b100011010;
				8'b1010001: c <= 9'b100111000;
				8'b1010100: c <= 9'b1111000;
				8'b1100110: c <= 9'b10100011;
				8'b101010: c <= 9'b11110110;
				8'b1011110: c <= 9'b100101110;
				8'b1100111: c <= 9'b10111;
				8'b1011010: c <= 9'b11001110;
				8'b1000010: c <= 9'b1110100;
				8'b111101: c <= 9'b111110011;
				8'b110000: c <= 9'b100110000;
				8'b111110: c <= 9'b1000011;
				8'b1100010: c <= 9'b101000101;
				8'b1110000: c <= 9'b111101100;
				8'b1101001: c <= 9'b10100011;
				8'b1110011: c <= 9'b101010000;
				8'b1001100: c <= 9'b100000011;
				8'b100001: c <= 9'b101101001;
				8'b1000110: c <= 9'b111011100;
				8'b1110010: c <= 9'b110010010;
				8'b1010000: c <= 9'b100110;
				8'b1111010: c <= 9'b110100001;
				8'b1010101: c <= 9'b101110110;
				8'b111011: c <= 9'b11011000;
				8'b1001101: c <= 9'b101101101;
				8'b111111: c <= 9'b100111001;
				8'b1101110: c <= 9'b101001100;
				8'b1111011: c <= 9'b101010010;
				8'b1001011: c <= 9'b101001000;
				8'b1101111: c <= 9'b100110100;
				8'b1101000: c <= 9'b111101100;
				8'b101100: c <= 9'b111001;
				8'b100100: c <= 9'b100;
				8'b1111000: c <= 9'b110101100;
				8'b1000101: c <= 9'b11100010;
				8'b1011001: c <= 9'b1101;
				8'b110100: c <= 9'b111011;
				8'b1111001: c <= 9'b10010110;
				8'b1110001: c <= 9'b1101010;
				8'b1001111: c <= 9'b111110101;
				8'b1100101: c <= 9'b11010100;
				8'b1111110: c <= 9'b100101000;
				8'b1111100: c <= 9'b1011110;
				8'b1010110: c <= 9'b110110100;
				8'b110010: c <= 9'b11010000;
				8'b1101101: c <= 9'b101110110;
				8'b100011: c <= 9'b11111001;
				8'b1110101: c <= 9'b110010110;
				8'b1111101: c <= 9'b101100110;
				8'b101001: c <= 9'b10001110;
				8'b1010010: c <= 9'b1011111;
				8'b1011000: c <= 9'b11111101;
				8'b101110: c <= 9'b110110010;
				8'b1000001: c <= 9'b11011000;
				default: c <= 9'b0;
			endcase
			9'b10000110 : case(di)
				8'b1000011: c <= 9'b11011010;
				8'b101000: c <= 9'b10110111;
				8'b111010: c <= 9'b111100011;
				8'b110110: c <= 9'b111010000;
				8'b1100100: c <= 9'b110101;
				8'b1000000: c <= 9'b10000101;
				8'b1110110: c <= 9'b1011111;
				8'b100101: c <= 9'b11000111;
				8'b101111: c <= 9'b10100101;
				8'b100110: c <= 9'b11111100;
				8'b1100011: c <= 9'b1111000;
				8'b1001000: c <= 9'b10101111;
				8'b111000: c <= 9'b11010;
				8'b110001: c <= 9'b11100111;
				8'b1010111: c <= 9'b110011000;
				8'b1001110: c <= 9'b1111011;
				8'b1101010: c <= 9'b111000;
				8'b1001001: c <= 9'b100010100;
				8'b1100000: c <= 9'b11000000;
				8'b110111: c <= 9'b100010010;
				8'b1011101: c <= 9'b111000110;
				8'b1011011: c <= 9'b100100001;
				8'b111001: c <= 9'b10000001;
				8'b1001010: c <= 9'b110000011;
				8'b110011: c <= 9'b1100001;
				8'b1101100: c <= 9'b100001110;
				8'b1110111: c <= 9'b100101001;
				8'b101011: c <= 9'b101110000;
				8'b1101011: c <= 9'b110001101;
				8'b111100: c <= 9'b10000111;
				8'b1000111: c <= 9'b111000101;
				8'b1011111: c <= 9'b100010110;
				8'b1110100: c <= 9'b110001101;
				8'b101101: c <= 9'b1100001;
				8'b1010011: c <= 9'b1101110;
				8'b1100001: c <= 9'b111001100;
				8'b110101: c <= 9'b100111000;
				8'b1000100: c <= 9'b11100011;
				8'b1010001: c <= 9'b101011111;
				8'b1010100: c <= 9'b110011011;
				8'b1100110: c <= 9'b110000;
				8'b101010: c <= 9'b11101100;
				8'b1011110: c <= 9'b1100010;
				8'b1100111: c <= 9'b10101;
				8'b1011010: c <= 9'b11110010;
				8'b1000010: c <= 9'b110001000;
				8'b111101: c <= 9'b1111000;
				8'b110000: c <= 9'b110111;
				8'b111110: c <= 9'b11001111;
				8'b1100010: c <= 9'b100110110;
				8'b1110000: c <= 9'b111001000;
				8'b1101001: c <= 9'b10101110;
				8'b1110011: c <= 9'b100111111;
				8'b1001100: c <= 9'b11010000;
				8'b100001: c <= 9'b110011;
				8'b1000110: c <= 9'b100101000;
				8'b1110010: c <= 9'b110101101;
				8'b1010000: c <= 9'b110110000;
				8'b1111010: c <= 9'b100001101;
				8'b1010101: c <= 9'b11011101;
				8'b111011: c <= 9'b101011000;
				8'b1001101: c <= 9'b111001000;
				8'b111111: c <= 9'b110011001;
				8'b1101110: c <= 9'b11100000;
				8'b1111011: c <= 9'b1100000;
				8'b1001011: c <= 9'b11011110;
				8'b1101111: c <= 9'b110110011;
				8'b1101000: c <= 9'b10110010;
				8'b101100: c <= 9'b111111110;
				8'b100100: c <= 9'b111101;
				8'b1111000: c <= 9'b11011011;
				8'b1000101: c <= 9'b10;
				8'b1011001: c <= 9'b111001010;
				8'b110100: c <= 9'b100011000;
				8'b1111001: c <= 9'b1100111;
				8'b1110001: c <= 9'b111110001;
				8'b1001111: c <= 9'b111100;
				8'b1100101: c <= 9'b100111110;
				8'b1111110: c <= 9'b10011111;
				8'b1111100: c <= 9'b10101011;
				8'b1010110: c <= 9'b11110100;
				8'b110010: c <= 9'b101110001;
				8'b1101101: c <= 9'b100101011;
				8'b100011: c <= 9'b110000010;
				8'b1110101: c <= 9'b11110100;
				8'b1111101: c <= 9'b100111000;
				8'b101001: c <= 9'b11110101;
				8'b1010010: c <= 9'b110110110;
				8'b1011000: c <= 9'b11000000;
				8'b101110: c <= 9'b100100010;
				8'b1000001: c <= 9'b101101;
				default: c <= 9'b0;
			endcase
			9'b10100010 : case(di)
				8'b1000011: c <= 9'b100001110;
				8'b101000: c <= 9'b10101000;
				8'b111010: c <= 9'b10011101;
				8'b110110: c <= 9'b10001110;
				8'b1100100: c <= 9'b10111;
				8'b1000000: c <= 9'b1001110;
				8'b1110110: c <= 9'b110111111;
				8'b100101: c <= 9'b1010000;
				8'b101111: c <= 9'b100110010;
				8'b100110: c <= 9'b110010011;
				8'b1100011: c <= 9'b100111001;
				8'b1001000: c <= 9'b100111;
				8'b111000: c <= 9'b111010010;
				8'b110001: c <= 9'b111011010;
				8'b1010111: c <= 9'b100010100;
				8'b1001110: c <= 9'b100111;
				8'b1101010: c <= 9'b100100000;
				8'b1001001: c <= 9'b100000110;
				8'b1100000: c <= 9'b100100010;
				8'b110111: c <= 9'b101000;
				8'b1011101: c <= 9'b111100011;
				8'b1011011: c <= 9'b10110011;
				8'b111001: c <= 9'b1000000;
				8'b1001010: c <= 9'b1001;
				8'b110011: c <= 9'b1101001;
				8'b1101100: c <= 9'b101100;
				8'b1110111: c <= 9'b100001100;
				8'b101011: c <= 9'b110100010;
				8'b1101011: c <= 9'b111000111;
				8'b111100: c <= 9'b11010000;
				8'b1000111: c <= 9'b100101011;
				8'b1011111: c <= 9'b11000100;
				8'b1110100: c <= 9'b111101110;
				8'b101101: c <= 9'b100011;
				8'b1010011: c <= 9'b100000100;
				8'b1100001: c <= 9'b110110110;
				8'b110101: c <= 9'b11000011;
				8'b1000100: c <= 9'b1100111;
				8'b1010001: c <= 9'b111001011;
				8'b1010100: c <= 9'b100001101;
				8'b1100110: c <= 9'b10111;
				8'b101010: c <= 9'b111101;
				8'b1011110: c <= 9'b101100100;
				8'b1100111: c <= 9'b110100;
				8'b1011010: c <= 9'b110010100;
				8'b1000010: c <= 9'b100011101;
				8'b111101: c <= 9'b101100000;
				8'b110000: c <= 9'b110010110;
				8'b111110: c <= 9'b1101101;
				8'b1100010: c <= 9'b110001011;
				8'b1110000: c <= 9'b10101011;
				8'b1101001: c <= 9'b111100101;
				8'b1110011: c <= 9'b100101010;
				8'b1001100: c <= 9'b110100110;
				8'b100001: c <= 9'b10111111;
				8'b1000110: c <= 9'b11011;
				8'b1110010: c <= 9'b100100011;
				8'b1010000: c <= 9'b100001101;
				8'b1111010: c <= 9'b10101000;
				8'b1010101: c <= 9'b1000;
				8'b111011: c <= 9'b100111110;
				8'b1001101: c <= 9'b110011100;
				8'b111111: c <= 9'b10011101;
				8'b1101110: c <= 9'b10000000;
				8'b1111011: c <= 9'b101110001;
				8'b1001011: c <= 9'b111010000;
				8'b1101111: c <= 9'b110101;
				8'b1101000: c <= 9'b10010000;
				8'b101100: c <= 9'b10101010;
				8'b100100: c <= 9'b10010110;
				8'b1111000: c <= 9'b100001010;
				8'b1000101: c <= 9'b100010011;
				8'b1011001: c <= 9'b110000;
				8'b110100: c <= 9'b100000110;
				8'b1111001: c <= 9'b11111010;
				8'b1110001: c <= 9'b11011;
				8'b1001111: c <= 9'b1001010;
				8'b1100101: c <= 9'b100100011;
				8'b1111110: c <= 9'b11110010;
				8'b1111100: c <= 9'b11100110;
				8'b1010110: c <= 9'b11000000;
				8'b110010: c <= 9'b11000110;
				8'b1101101: c <= 9'b11001101;
				8'b100011: c <= 9'b110111;
				8'b1110101: c <= 9'b110010011;
				8'b1111101: c <= 9'b101110011;
				8'b101001: c <= 9'b11010;
				8'b1010010: c <= 9'b1000001;
				8'b1011000: c <= 9'b100000101;
				8'b101110: c <= 9'b100010;
				8'b1000001: c <= 9'b111111;
				default: c <= 9'b0;
			endcase
			9'b101111001 : case(di)
				8'b1000011: c <= 9'b110110111;
				8'b101000: c <= 9'b101010000;
				8'b111010: c <= 9'b111101101;
				8'b110110: c <= 9'b11101000;
				8'b1100100: c <= 9'b101101100;
				8'b1000000: c <= 9'b111001001;
				8'b1110110: c <= 9'b101110110;
				8'b100101: c <= 9'b100101000;
				8'b101111: c <= 9'b111100011;
				8'b100110: c <= 9'b111010;
				8'b1100011: c <= 9'b111101010;
				8'b1001000: c <= 9'b10000101;
				8'b111000: c <= 9'b1001110;
				8'b110001: c <= 9'b10010111;
				8'b1010111: c <= 9'b10010011;
				8'b1001110: c <= 9'b100001100;
				8'b1101010: c <= 9'b100011101;
				8'b1001001: c <= 9'b110101;
				8'b1100000: c <= 9'b101000110;
				8'b110111: c <= 9'b101001110;
				8'b1011101: c <= 9'b111011;
				8'b1011011: c <= 9'b11111010;
				8'b111001: c <= 9'b11001000;
				8'b1001010: c <= 9'b111001100;
				8'b110011: c <= 9'b11000010;
				8'b1101100: c <= 9'b111010010;
				8'b1110111: c <= 9'b101101000;
				8'b101011: c <= 9'b110110010;
				8'b1101011: c <= 9'b10011100;
				8'b111100: c <= 9'b10110010;
				8'b1000111: c <= 9'b100110111;
				8'b1011111: c <= 9'b10000110;
				8'b1110100: c <= 9'b111011111;
				8'b101101: c <= 9'b111001010;
				8'b1010011: c <= 9'b110101001;
				8'b1100001: c <= 9'b11100101;
				8'b110101: c <= 9'b1100110;
				8'b1000100: c <= 9'b11110000;
				8'b1010001: c <= 9'b111101;
				8'b1010100: c <= 9'b1011100;
				8'b1100110: c <= 9'b110010;
				8'b101010: c <= 9'b110010111;
				8'b1011110: c <= 9'b110111011;
				8'b1100111: c <= 9'b101000001;
				8'b1011010: c <= 9'b110100010;
				8'b1000010: c <= 9'b101110101;
				8'b111101: c <= 9'b101100111;
				8'b110000: c <= 9'b11000110;
				8'b111110: c <= 9'b101011101;
				8'b1100010: c <= 9'b100010111;
				8'b1110000: c <= 9'b10011100;
				8'b1101001: c <= 9'b101010101;
				8'b1110011: c <= 9'b110010010;
				8'b1001100: c <= 9'b1111110;
				8'b100001: c <= 9'b10000011;
				8'b1000110: c <= 9'b100001010;
				8'b1110010: c <= 9'b110010011;
				8'b1010000: c <= 9'b101011010;
				8'b1111010: c <= 9'b11;
				8'b1010101: c <= 9'b101011;
				8'b111011: c <= 9'b111000110;
				8'b1001101: c <= 9'b110111011;
				8'b111111: c <= 9'b1011000;
				8'b1101110: c <= 9'b100111001;
				8'b1111011: c <= 9'b111000010;
				8'b1001011: c <= 9'b11101101;
				8'b1101111: c <= 9'b111010111;
				8'b1101000: c <= 9'b100010101;
				8'b101100: c <= 9'b1010111;
				8'b100100: c <= 9'b111111101;
				8'b1111000: c <= 9'b10010;
				8'b1000101: c <= 9'b100110111;
				8'b1011001: c <= 9'b11010;
				8'b110100: c <= 9'b110100011;
				8'b1111001: c <= 9'b10101100;
				8'b1110001: c <= 9'b11011001;
				8'b1001111: c <= 9'b10011001;
				8'b1100101: c <= 9'b1111110;
				8'b1111110: c <= 9'b100011000;
				8'b1111100: c <= 9'b100111;
				8'b1010110: c <= 9'b100010001;
				8'b110010: c <= 9'b11000001;
				8'b1101101: c <= 9'b101000101;
				8'b100011: c <= 9'b1010000;
				8'b1110101: c <= 9'b110;
				8'b1111101: c <= 9'b10011000;
				8'b101001: c <= 9'b111110101;
				8'b1010010: c <= 9'b100110;
				8'b1011000: c <= 9'b100011101;
				8'b101110: c <= 9'b1001111;
				8'b1000001: c <= 9'b1110101;
				default: c <= 9'b0;
			endcase
			9'b111011 : case(di)
				8'b1000011: c <= 9'b101010;
				8'b101000: c <= 9'b10110001;
				8'b111010: c <= 9'b110111011;
				8'b110110: c <= 9'b1001001;
				8'b1100100: c <= 9'b10001010;
				8'b1000000: c <= 9'b101100000;
				8'b1110110: c <= 9'b11000000;
				8'b100101: c <= 9'b111110101;
				8'b101111: c <= 9'b110100100;
				8'b100110: c <= 9'b100010;
				8'b1100011: c <= 9'b101001100;
				8'b1001000: c <= 9'b1110111;
				8'b111000: c <= 9'b100000101;
				8'b110001: c <= 9'b11111;
				8'b1010111: c <= 9'b111001110;
				8'b1001110: c <= 9'b10101000;
				8'b1101010: c <= 9'b10111100;
				8'b1001001: c <= 9'b100010110;
				8'b1100000: c <= 9'b101000110;
				8'b110111: c <= 9'b10101;
				8'b1011101: c <= 9'b100101000;
				8'b1011011: c <= 9'b1000011;
				8'b111001: c <= 9'b110000011;
				8'b1001010: c <= 9'b1100111;
				8'b110011: c <= 9'b10;
				8'b1101100: c <= 9'b1001001;
				8'b1110111: c <= 9'b1010010;
				8'b101011: c <= 9'b1101100;
				8'b1101011: c <= 9'b110001011;
				8'b111100: c <= 9'b111011010;
				8'b1000111: c <= 9'b110101111;
				8'b1011111: c <= 9'b100101111;
				8'b1110100: c <= 9'b110000101;
				8'b101101: c <= 9'b100000100;
				8'b1010011: c <= 9'b1100111;
				8'b1100001: c <= 9'b101101;
				8'b110101: c <= 9'b100101;
				8'b1000100: c <= 9'b10011011;
				8'b1010001: c <= 9'b100101100;
				8'b1010100: c <= 9'b10000000;
				8'b1100110: c <= 9'b1;
				8'b101010: c <= 9'b10111100;
				8'b1011110: c <= 9'b10111100;
				8'b1100111: c <= 9'b10110;
				8'b1011010: c <= 9'b101010101;
				8'b1000010: c <= 9'b100001110;
				8'b111101: c <= 9'b11010001;
				8'b110000: c <= 9'b101000100;
				8'b111110: c <= 9'b10101010;
				8'b1100010: c <= 9'b110000011;
				8'b1110000: c <= 9'b10101111;
				8'b1101001: c <= 9'b11100110;
				8'b1110011: c <= 9'b10011;
				8'b1001100: c <= 9'b100000101;
				8'b100001: c <= 9'b110101110;
				8'b1000110: c <= 9'b101011010;
				8'b1110010: c <= 9'b111001011;
				8'b1010000: c <= 9'b1011111;
				8'b1111010: c <= 9'b110110111;
				8'b1010101: c <= 9'b10111011;
				8'b111011: c <= 9'b100101011;
				8'b1001101: c <= 9'b111001010;
				8'b111111: c <= 9'b100001011;
				8'b1101110: c <= 9'b110011001;
				8'b1111011: c <= 9'b101000101;
				8'b1001011: c <= 9'b11000011;
				8'b1101111: c <= 9'b11001100;
				8'b1101000: c <= 9'b111110110;
				8'b101100: c <= 9'b111000011;
				8'b100100: c <= 9'b1001101;
				8'b1111000: c <= 9'b100111010;
				8'b1000101: c <= 9'b101110001;
				8'b1011001: c <= 9'b100011;
				8'b110100: c <= 9'b101101001;
				8'b1111001: c <= 9'b10101110;
				8'b1110001: c <= 9'b111000010;
				8'b1001111: c <= 9'b1110101;
				8'b1100101: c <= 9'b111111000;
				8'b1111110: c <= 9'b100001100;
				8'b1111100: c <= 9'b10011010;
				8'b1010110: c <= 9'b111111000;
				8'b110010: c <= 9'b100001;
				8'b1101101: c <= 9'b101000101;
				8'b100011: c <= 9'b1001100;
				8'b1110101: c <= 9'b10100101;
				8'b1111101: c <= 9'b111100111;
				8'b101001: c <= 9'b11011000;
				8'b1010010: c <= 9'b1101111;
				8'b1011000: c <= 9'b100001;
				8'b101110: c <= 9'b100011011;
				8'b1000001: c <= 9'b101100001;
				default: c <= 9'b0;
			endcase
			9'b100111001 : case(di)
				8'b1000011: c <= 9'b100000010;
				8'b101000: c <= 9'b100001110;
				8'b111010: c <= 9'b100011;
				8'b110110: c <= 9'b100011000;
				8'b1100100: c <= 9'b11010100;
				8'b1000000: c <= 9'b110000000;
				8'b1110110: c <= 9'b110100111;
				8'b100101: c <= 9'b101110110;
				8'b101111: c <= 9'b100010001;
				8'b100110: c <= 9'b101000100;
				8'b1100011: c <= 9'b1;
				8'b1001000: c <= 9'b100000000;
				8'b111000: c <= 9'b1000100;
				8'b110001: c <= 9'b1000000;
				8'b1010111: c <= 9'b1101;
				8'b1001110: c <= 9'b100010010;
				8'b1101010: c <= 9'b110100011;
				8'b1001001: c <= 9'b100100010;
				8'b1100000: c <= 9'b1110000;
				8'b110111: c <= 9'b101010110;
				8'b1011101: c <= 9'b110100001;
				8'b1011011: c <= 9'b100000110;
				8'b111001: c <= 9'b110010110;
				8'b1001010: c <= 9'b100001001;
				8'b110011: c <= 9'b11100000;
				8'b1101100: c <= 9'b10101010;
				8'b1110111: c <= 9'b110001011;
				8'b101011: c <= 9'b111110011;
				8'b1101011: c <= 9'b101100010;
				8'b111100: c <= 9'b101001;
				8'b1000111: c <= 9'b10100101;
				8'b1011111: c <= 9'b1010010;
				8'b1110100: c <= 9'b11010011;
				8'b101101: c <= 9'b1001010;
				8'b1010011: c <= 9'b10110010;
				8'b1100001: c <= 9'b11011001;
				8'b110101: c <= 9'b11001000;
				8'b1000100: c <= 9'b110100000;
				8'b1010001: c <= 9'b1101101;
				8'b1010100: c <= 9'b11100111;
				8'b1100110: c <= 9'b110111011;
				8'b101010: c <= 9'b11001;
				8'b1011110: c <= 9'b101101;
				8'b1100111: c <= 9'b101011110;
				8'b1011010: c <= 9'b10000011;
				8'b1000010: c <= 9'b101010101;
				8'b111101: c <= 9'b100000111;
				8'b110000: c <= 9'b110001100;
				8'b111110: c <= 9'b10110110;
				8'b1100010: c <= 9'b111111110;
				8'b1110000: c <= 9'b10010111;
				8'b1101001: c <= 9'b101111110;
				8'b1110011: c <= 9'b101100001;
				8'b1001100: c <= 9'b101100111;
				8'b100001: c <= 9'b11011;
				8'b1000110: c <= 9'b10111011;
				8'b1110010: c <= 9'b10011100;
				8'b1010000: c <= 9'b101010011;
				8'b1111010: c <= 9'b110101110;
				8'b1010101: c <= 9'b110101001;
				8'b111011: c <= 9'b100000011;
				8'b1001101: c <= 9'b1011011;
				8'b111111: c <= 9'b110110101;
				8'b1101110: c <= 9'b100001101;
				8'b1111011: c <= 9'b100010101;
				8'b1001011: c <= 9'b110000101;
				8'b1101111: c <= 9'b110101010;
				8'b1101000: c <= 9'b1101110;
				8'b101100: c <= 9'b111011111;
				8'b100100: c <= 9'b11111101;
				8'b1111000: c <= 9'b110010011;
				8'b1000101: c <= 9'b110100;
				8'b1011001: c <= 9'b110000001;
				8'b110100: c <= 9'b100111010;
				8'b1111001: c <= 9'b11101111;
				8'b1110001: c <= 9'b101011000;
				8'b1001111: c <= 9'b11010;
				8'b1100101: c <= 9'b101010111;
				8'b1111110: c <= 9'b111011111;
				8'b1111100: c <= 9'b111001011;
				8'b1010110: c <= 9'b100111001;
				8'b110010: c <= 9'b11;
				8'b1101101: c <= 9'b111001010;
				8'b100011: c <= 9'b111101001;
				8'b1110101: c <= 9'b1111;
				8'b1111101: c <= 9'b101110110;
				8'b101001: c <= 9'b101000111;
				8'b1010010: c <= 9'b110101010;
				8'b1011000: c <= 9'b11101000;
				8'b101110: c <= 9'b10000011;
				8'b1000001: c <= 9'b101100;
				default: c <= 9'b0;
			endcase
			9'b11111011 : case(di)
				8'b1000011: c <= 9'b100111000;
				8'b101000: c <= 9'b10100011;
				8'b111010: c <= 9'b100010011;
				8'b110110: c <= 9'b10101011;
				8'b1100100: c <= 9'b101100101;
				8'b1000000: c <= 9'b1001011;
				8'b1110110: c <= 9'b101010000;
				8'b100101: c <= 9'b110001101;
				8'b101111: c <= 9'b1001;
				8'b100110: c <= 9'b101001000;
				8'b1100011: c <= 9'b101011000;
				8'b1001000: c <= 9'b101011101;
				8'b111000: c <= 9'b101100010;
				8'b110001: c <= 9'b101110110;
				8'b1010111: c <= 9'b110100001;
				8'b1001110: c <= 9'b1100;
				8'b1101010: c <= 9'b101111110;
				8'b1001001: c <= 9'b10000101;
				8'b1100000: c <= 9'b111110011;
				8'b110111: c <= 9'b110000111;
				8'b1011101: c <= 9'b110100101;
				8'b1011011: c <= 9'b11111000;
				8'b111001: c <= 9'b10011111;
				8'b1001010: c <= 9'b100111100;
				8'b110011: c <= 9'b10100110;
				8'b1101100: c <= 9'b10010101;
				8'b1110111: c <= 9'b11100000;
				8'b101011: c <= 9'b110111;
				8'b1101011: c <= 9'b1001011;
				8'b111100: c <= 9'b1010011;
				8'b1000111: c <= 9'b100100001;
				8'b1011111: c <= 9'b11001100;
				8'b1110100: c <= 9'b11010011;
				8'b101101: c <= 9'b101100010;
				8'b1010011: c <= 9'b1000001;
				8'b1100001: c <= 9'b100101010;
				8'b110101: c <= 9'b1110001;
				8'b1000100: c <= 9'b11010011;
				8'b1010001: c <= 9'b101101011;
				8'b1010100: c <= 9'b11001010;
				8'b1100110: c <= 9'b10000011;
				8'b101010: c <= 9'b10111;
				8'b1011110: c <= 9'b10011101;
				8'b1100111: c <= 9'b10100101;
				8'b1011010: c <= 9'b111010001;
				8'b1000010: c <= 9'b10;
				8'b111101: c <= 9'b11101001;
				8'b110000: c <= 9'b111000110;
				8'b111110: c <= 9'b11101000;
				8'b1100010: c <= 9'b10111001;
				8'b1110000: c <= 9'b101111000;
				8'b1101001: c <= 9'b100010001;
				8'b1110011: c <= 9'b11100111;
				8'b1001100: c <= 9'b11011110;
				8'b100001: c <= 9'b101100011;
				8'b1000110: c <= 9'b11110;
				8'b1110010: c <= 9'b101001111;
				8'b1010000: c <= 9'b111101111;
				8'b1111010: c <= 9'b111101101;
				8'b1010101: c <= 9'b101100011;
				8'b111011: c <= 9'b100010110;
				8'b1001101: c <= 9'b10;
				8'b111111: c <= 9'b100000010;
				8'b1101110: c <= 9'b111100110;
				8'b1111011: c <= 9'b101000010;
				8'b1001011: c <= 9'b11011110;
				8'b1101111: c <= 9'b10110;
				8'b1101000: c <= 9'b11001101;
				8'b101100: c <= 9'b11011010;
				8'b100100: c <= 9'b111101000;
				8'b1111000: c <= 9'b101011;
				8'b1000101: c <= 9'b1101;
				8'b1011001: c <= 9'b101010110;
				8'b110100: c <= 9'b11011000;
				8'b1111001: c <= 9'b111110110;
				8'b1110001: c <= 9'b11011;
				8'b1001111: c <= 9'b1000000;
				8'b1100101: c <= 9'b100001110;
				8'b1111110: c <= 9'b11011101;
				8'b1111100: c <= 9'b10100000;
				8'b1010110: c <= 9'b101010011;
				8'b110010: c <= 9'b101010010;
				8'b1101101: c <= 9'b100101111;
				8'b100011: c <= 9'b101101011;
				8'b1110101: c <= 9'b10111;
				8'b1111101: c <= 9'b1010010;
				8'b101001: c <= 9'b1101100;
				8'b1010010: c <= 9'b111011010;
				8'b1011000: c <= 9'b10011010;
				8'b101110: c <= 9'b110100001;
				8'b1000001: c <= 9'b101001111;
				default: c <= 9'b0;
			endcase
			9'b1011100 : case(di)
				8'b1000011: c <= 9'b10000110;
				8'b101000: c <= 9'b1101010;
				8'b111010: c <= 9'b10101;
				8'b110110: c <= 9'b111011101;
				8'b1100100: c <= 9'b1101000;
				8'b1000000: c <= 9'b100000011;
				8'b1110110: c <= 9'b11110100;
				8'b100101: c <= 9'b100000110;
				8'b101111: c <= 9'b11100010;
				8'b100110: c <= 9'b1010010;
				8'b1100011: c <= 9'b11111;
				8'b1001000: c <= 9'b110100101;
				8'b111000: c <= 9'b11010000;
				8'b110001: c <= 9'b101010000;
				8'b1010111: c <= 9'b1011011;
				8'b1001110: c <= 9'b11111110;
				8'b1101010: c <= 9'b1101100;
				8'b1001001: c <= 9'b1100101;
				8'b1100000: c <= 9'b110010001;
				8'b110111: c <= 9'b111010001;
				8'b1011101: c <= 9'b11110010;
				8'b1011011: c <= 9'b111000000;
				8'b111001: c <= 9'b11111011;
				8'b1001010: c <= 9'b111101001;
				8'b110011: c <= 9'b101010101;
				8'b1101100: c <= 9'b111000000;
				8'b1110111: c <= 9'b1101101;
				8'b101011: c <= 9'b10000110;
				8'b1101011: c <= 9'b100001100;
				8'b111100: c <= 9'b111011011;
				8'b1000111: c <= 9'b10010101;
				8'b1011111: c <= 9'b100000111;
				8'b1110100: c <= 9'b111100011;
				8'b101101: c <= 9'b100001;
				8'b1010011: c <= 9'b111100101;
				8'b1100001: c <= 9'b111100110;
				8'b110101: c <= 9'b101001110;
				8'b1000100: c <= 9'b100000010;
				8'b1010001: c <= 9'b11001110;
				8'b1010100: c <= 9'b101;
				8'b1100110: c <= 9'b101101000;
				8'b101010: c <= 9'b111010;
				8'b1011110: c <= 9'b11111001;
				8'b1100111: c <= 9'b101000100;
				8'b1011010: c <= 9'b110011010;
				8'b1000010: c <= 9'b100101110;
				8'b111101: c <= 9'b1101010;
				8'b110000: c <= 9'b10000011;
				8'b111110: c <= 9'b100011010;
				8'b1100010: c <= 9'b11100100;
				8'b1110000: c <= 9'b111010110;
				8'b1101001: c <= 9'b101101110;
				8'b1110011: c <= 9'b100010000;
				8'b1001100: c <= 9'b100001001;
				8'b100001: c <= 9'b100100101;
				8'b1000110: c <= 9'b111011110;
				8'b1110010: c <= 9'b111011;
				8'b1010000: c <= 9'b110011111;
				8'b1111010: c <= 9'b1001000;
				8'b1010101: c <= 9'b10101101;
				8'b111011: c <= 9'b111010100;
				8'b1001101: c <= 9'b100000110;
				8'b111111: c <= 9'b10010101;
				8'b1101110: c <= 9'b110111011;
				8'b1111011: c <= 9'b11011110;
				8'b1001011: c <= 9'b1111000;
				8'b1101111: c <= 9'b100100000;
				8'b1101000: c <= 9'b10001000;
				8'b101100: c <= 9'b110101010;
				8'b100100: c <= 9'b10110111;
				8'b1111000: c <= 9'b101011010;
				8'b1000101: c <= 9'b110100001;
				8'b1011001: c <= 9'b10100;
				8'b110100: c <= 9'b11101101;
				8'b1111001: c <= 9'b100111011;
				8'b1110001: c <= 9'b111110110;
				8'b1001111: c <= 9'b111000101;
				8'b1100101: c <= 9'b100110101;
				8'b1111110: c <= 9'b100001001;
				8'b1111100: c <= 9'b110100;
				8'b1010110: c <= 9'b10101;
				8'b110010: c <= 9'b100100110;
				8'b1101101: c <= 9'b100110111;
				8'b100011: c <= 9'b100110111;
				8'b1110101: c <= 9'b11110101;
				8'b1111101: c <= 9'b111000010;
				8'b101001: c <= 9'b100010110;
				8'b1010010: c <= 9'b11111;
				8'b1011000: c <= 9'b1111101;
				8'b101110: c <= 9'b11011101;
				8'b1000001: c <= 9'b110000000;
				default: c <= 9'b0;
			endcase
			9'b110000110 : case(di)
				8'b1000011: c <= 9'b1010011;
				8'b101000: c <= 9'b101011101;
				8'b111010: c <= 9'b11001001;
				8'b110110: c <= 9'b101000010;
				8'b1100100: c <= 9'b101101100;
				8'b1000000: c <= 9'b111100001;
				8'b1110110: c <= 9'b100111111;
				8'b100101: c <= 9'b10101100;
				8'b101111: c <= 9'b10101010;
				8'b100110: c <= 9'b101001000;
				8'b1100011: c <= 9'b101010111;
				8'b1001000: c <= 9'b100010000;
				8'b111000: c <= 9'b101101011;
				8'b110001: c <= 9'b10011100;
				8'b1010111: c <= 9'b111100101;
				8'b1001110: c <= 9'b110101111;
				8'b1101010: c <= 9'b101010000;
				8'b1001001: c <= 9'b101101001;
				8'b1100000: c <= 9'b100111110;
				8'b110111: c <= 9'b101001000;
				8'b1011101: c <= 9'b100;
				8'b1011011: c <= 9'b100001110;
				8'b111001: c <= 9'b101010100;
				8'b1001010: c <= 9'b100011101;
				8'b110011: c <= 9'b11000;
				8'b1101100: c <= 9'b101001100;
				8'b1110111: c <= 9'b10001110;
				8'b101011: c <= 9'b111101010;
				8'b1101011: c <= 9'b101010011;
				8'b111100: c <= 9'b10101010;
				8'b1000111: c <= 9'b1001011;
				8'b1011111: c <= 9'b11010011;
				8'b1110100: c <= 9'b100110;
				8'b101101: c <= 9'b1011;
				8'b1010011: c <= 9'b100011111;
				8'b1100001: c <= 9'b101110110;
				8'b110101: c <= 9'b100001111;
				8'b1000100: c <= 9'b10010111;
				8'b1010001: c <= 9'b11111000;
				8'b1010100: c <= 9'b1100111;
				8'b1100110: c <= 9'b1111001;
				8'b101010: c <= 9'b1011;
				8'b1011110: c <= 9'b10110001;
				8'b1100111: c <= 9'b100011;
				8'b1011010: c <= 9'b1000000;
				8'b1000010: c <= 9'b110000010;
				8'b111101: c <= 9'b10101100;
				8'b110000: c <= 9'b11100;
				8'b111110: c <= 9'b11000110;
				8'b1100010: c <= 9'b100011100;
				8'b1110000: c <= 9'b10110100;
				8'b1101001: c <= 9'b11000110;
				8'b1110011: c <= 9'b1110100;
				8'b1001100: c <= 9'b101011110;
				8'b100001: c <= 9'b11110001;
				8'b1000110: c <= 9'b1110100;
				8'b1110010: c <= 9'b110011;
				8'b1010000: c <= 9'b1011001;
				8'b1111010: c <= 9'b1011010;
				8'b1010101: c <= 9'b110011001;
				8'b111011: c <= 9'b111000;
				8'b1001101: c <= 9'b111101100;
				8'b111111: c <= 9'b100101000;
				8'b1101110: c <= 9'b111010111;
				8'b1111011: c <= 9'b11000001;
				8'b1001011: c <= 9'b100001010;
				8'b1101111: c <= 9'b1100000;
				8'b1101000: c <= 9'b111111;
				8'b101100: c <= 9'b11111100;
				8'b100100: c <= 9'b11110011;
				8'b1111000: c <= 9'b110100111;
				8'b1000101: c <= 9'b1010010;
				8'b1011001: c <= 9'b101100100;
				8'b110100: c <= 9'b111011100;
				8'b1111001: c <= 9'b101010000;
				8'b1110001: c <= 9'b101000011;
				8'b1001111: c <= 9'b1111010;
				8'b1100101: c <= 9'b1011001;
				8'b1111110: c <= 9'b11100010;
				8'b1111100: c <= 9'b1101;
				8'b1010110: c <= 9'b11101101;
				8'b110010: c <= 9'b10101011;
				8'b1101101: c <= 9'b11011010;
				8'b100011: c <= 9'b110011011;
				8'b1110101: c <= 9'b100010100;
				8'b1111101: c <= 9'b1001100;
				8'b101001: c <= 9'b111000010;
				8'b1010010: c <= 9'b111111;
				8'b1011000: c <= 9'b111001001;
				8'b101110: c <= 9'b101101100;
				8'b1000001: c <= 9'b100100;
				default: c <= 9'b0;
			endcase
			9'b100100011 : case(di)
				8'b1000011: c <= 9'b11110001;
				8'b101000: c <= 9'b10110011;
				8'b111010: c <= 9'b1111010;
				8'b110110: c <= 9'b1;
				8'b1100100: c <= 9'b100100111;
				8'b1000000: c <= 9'b111100;
				8'b1110110: c <= 9'b100100101;
				8'b100101: c <= 9'b110100101;
				8'b101111: c <= 9'b110011001;
				8'b100110: c <= 9'b110011000;
				8'b1100011: c <= 9'b11010000;
				8'b1001000: c <= 9'b1011011;
				8'b111000: c <= 9'b111101111;
				8'b110001: c <= 9'b1101110;
				8'b1010111: c <= 9'b111010111;
				8'b1001110: c <= 9'b111010111;
				8'b1101010: c <= 9'b101011101;
				8'b1001001: c <= 9'b111001011;
				8'b1100000: c <= 9'b11011100;
				8'b110111: c <= 9'b11111100;
				8'b1011101: c <= 9'b11110110;
				8'b1011011: c <= 9'b111010100;
				8'b111001: c <= 9'b1010111;
				8'b1001010: c <= 9'b1010011;
				8'b110011: c <= 9'b1011;
				8'b1101100: c <= 9'b100001001;
				8'b1110111: c <= 9'b110100001;
				8'b101011: c <= 9'b101100;
				8'b1101011: c <= 9'b10100110;
				8'b111100: c <= 9'b100000011;
				8'b1000111: c <= 9'b11111000;
				8'b1011111: c <= 9'b1001000;
				8'b1110100: c <= 9'b111110110;
				8'b101101: c <= 9'b1000001;
				8'b1010011: c <= 9'b1110111;
				8'b1100001: c <= 9'b111111010;
				8'b110101: c <= 9'b10110100;
				8'b1000100: c <= 9'b110001001;
				8'b1010001: c <= 9'b110110111;
				8'b1010100: c <= 9'b10110001;
				8'b1100110: c <= 9'b100110110;
				8'b101010: c <= 9'b1000100;
				8'b1011110: c <= 9'b110010011;
				8'b1100111: c <= 9'b100001111;
				8'b1011010: c <= 9'b111000000;
				8'b1000010: c <= 9'b10101;
				8'b111101: c <= 9'b10010100;
				8'b110000: c <= 9'b100001011;
				8'b111110: c <= 9'b111100000;
				8'b1100010: c <= 9'b111101111;
				8'b1110000: c <= 9'b111001101;
				8'b1101001: c <= 9'b100001101;
				8'b1110011: c <= 9'b110011111;
				8'b1001100: c <= 9'b100011;
				8'b100001: c <= 9'b101111000;
				8'b1000110: c <= 9'b110010101;
				8'b1110010: c <= 9'b1000001;
				8'b1010000: c <= 9'b101011101;
				8'b1111010: c <= 9'b100110111;
				8'b1010101: c <= 9'b100000011;
				8'b111011: c <= 9'b1001110;
				8'b1001101: c <= 9'b111100000;
				8'b111111: c <= 9'b11001100;
				8'b1101110: c <= 9'b11000;
				8'b1111011: c <= 9'b100001010;
				8'b1001011: c <= 9'b10100111;
				8'b1101111: c <= 9'b11111011;
				8'b1101000: c <= 9'b101110101;
				8'b101100: c <= 9'b111001001;
				8'b100100: c <= 9'b100011001;
				8'b1111000: c <= 9'b111100110;
				8'b1000101: c <= 9'b110110101;
				8'b1011001: c <= 9'b110010110;
				8'b110100: c <= 9'b110100111;
				8'b1111001: c <= 9'b11011001;
				8'b1110001: c <= 9'b1010010;
				8'b1001111: c <= 9'b10010111;
				8'b1100101: c <= 9'b100000110;
				8'b1111110: c <= 9'b111000111;
				8'b1111100: c <= 9'b1110010;
				8'b1010110: c <= 9'b101111001;
				8'b110010: c <= 9'b101011111;
				8'b1101101: c <= 9'b11001;
				8'b100011: c <= 9'b100101011;
				8'b1110101: c <= 9'b1101101;
				8'b1111101: c <= 9'b101100011;
				8'b101001: c <= 9'b100011111;
				8'b1010010: c <= 9'b101110101;
				8'b1011000: c <= 9'b110010100;
				8'b101110: c <= 9'b1000001;
				8'b1000001: c <= 9'b110000000;
				default: c <= 9'b0;
			endcase
			9'b1100100 : case(di)
				8'b1000011: c <= 9'b101101001;
				8'b101000: c <= 9'b101111110;
				8'b111010: c <= 9'b101010010;
				8'b110110: c <= 9'b110000011;
				8'b1100100: c <= 9'b100111001;
				8'b1000000: c <= 9'b10111010;
				8'b1110110: c <= 9'b111100101;
				8'b100101: c <= 9'b11110001;
				8'b101111: c <= 9'b1100011;
				8'b100110: c <= 9'b1100100;
				8'b1100011: c <= 9'b1111101;
				8'b1001000: c <= 9'b111011111;
				8'b111000: c <= 9'b111101111;
				8'b110001: c <= 9'b111001110;
				8'b1010111: c <= 9'b1110101;
				8'b1001110: c <= 9'b1111000;
				8'b1101010: c <= 9'b11001;
				8'b1001001: c <= 9'b10111000;
				8'b1100000: c <= 9'b111100010;
				8'b110111: c <= 9'b101001001;
				8'b1011101: c <= 9'b111001100;
				8'b1011011: c <= 9'b110101;
				8'b111001: c <= 9'b111101000;
				8'b1001010: c <= 9'b10010011;
				8'b110011: c <= 9'b101010111;
				8'b1101100: c <= 9'b10100110;
				8'b1110111: c <= 9'b11100010;
				8'b101011: c <= 9'b101001111;
				8'b1101011: c <= 9'b100001;
				8'b111100: c <= 9'b111011111;
				8'b1000111: c <= 9'b11111101;
				8'b1011111: c <= 9'b100111111;
				8'b1110100: c <= 9'b11110110;
				8'b101101: c <= 9'b111001010;
				8'b1010011: c <= 9'b100001;
				8'b1100001: c <= 9'b100010001;
				8'b110101: c <= 9'b100111101;
				8'b1000100: c <= 9'b11001000;
				8'b1010001: c <= 9'b110011011;
				8'b1010100: c <= 9'b110111010;
				8'b1100110: c <= 9'b1011111;
				8'b101010: c <= 9'b100110101;
				8'b1011110: c <= 9'b110001110;
				8'b1100111: c <= 9'b11101;
				8'b1011010: c <= 9'b111100110;
				8'b1000010: c <= 9'b10101;
				8'b111101: c <= 9'b100100010;
				8'b110000: c <= 9'b10111011;
				8'b111110: c <= 9'b1100010;
				8'b1100010: c <= 9'b110011;
				8'b1110000: c <= 9'b1000101;
				8'b1101001: c <= 9'b10010101;
				8'b1110011: c <= 9'b10001100;
				8'b1001100: c <= 9'b101011;
				8'b100001: c <= 9'b100110110;
				8'b1000110: c <= 9'b111110101;
				8'b1110010: c <= 9'b10101100;
				8'b1010000: c <= 9'b101101010;
				8'b1111010: c <= 9'b110101011;
				8'b1010101: c <= 9'b101000;
				8'b111011: c <= 9'b1011110;
				8'b1001101: c <= 9'b100110011;
				8'b111111: c <= 9'b111011100;
				8'b1101110: c <= 9'b11000011;
				8'b1111011: c <= 9'b11100110;
				8'b1001011: c <= 9'b110001001;
				8'b1101111: c <= 9'b11111010;
				8'b1101000: c <= 9'b110010100;
				8'b101100: c <= 9'b100111110;
				8'b100100: c <= 9'b101101010;
				8'b1111000: c <= 9'b11011000;
				8'b1000101: c <= 9'b101000010;
				8'b1011001: c <= 9'b1100010;
				8'b110100: c <= 9'b1001100;
				8'b1111001: c <= 9'b100011010;
				8'b1110001: c <= 9'b1100111;
				8'b1001111: c <= 9'b10001100;
				8'b1100101: c <= 9'b11101100;
				8'b1111110: c <= 9'b111010100;
				8'b1111100: c <= 9'b111011110;
				8'b1010110: c <= 9'b100001;
				8'b110010: c <= 9'b10001000;
				8'b1101101: c <= 9'b111111010;
				8'b100011: c <= 9'b100011010;
				8'b1110101: c <= 9'b10101110;
				8'b1111101: c <= 9'b101100110;
				8'b101001: c <= 9'b11101100;
				8'b1010010: c <= 9'b101000011;
				8'b1011000: c <= 9'b111111010;
				8'b101110: c <= 9'b111100000;
				8'b1000001: c <= 9'b11001100;
				default: c <= 9'b0;
			endcase
			9'b100111 : case(di)
				8'b1000011: c <= 9'b11011001;
				8'b101000: c <= 9'b1010110;
				8'b111010: c <= 9'b11010001;
				8'b110110: c <= 9'b101011101;
				8'b1100100: c <= 9'b110101010;
				8'b1000000: c <= 9'b110101110;
				8'b1110110: c <= 9'b1000111;
				8'b100101: c <= 9'b11001;
				8'b101111: c <= 9'b100001011;
				8'b100110: c <= 9'b100001111;
				8'b1100011: c <= 9'b1110001;
				8'b1001000: c <= 9'b1100011;
				8'b111000: c <= 9'b1010000;
				8'b110001: c <= 9'b11110111;
				8'b1010111: c <= 9'b10111000;
				8'b1001110: c <= 9'b11000110;
				8'b1101010: c <= 9'b10111001;
				8'b1001001: c <= 9'b101111000;
				8'b1100000: c <= 9'b10010101;
				8'b110111: c <= 9'b100111;
				8'b1011101: c <= 9'b100110010;
				8'b1011011: c <= 9'b1101110;
				8'b111001: c <= 9'b10101011;
				8'b1001010: c <= 9'b111110110;
				8'b110011: c <= 9'b111111001;
				8'b1101100: c <= 9'b1001100;
				8'b1110111: c <= 9'b11100101;
				8'b101011: c <= 9'b1001100;
				8'b1101011: c <= 9'b110000010;
				8'b111100: c <= 9'b11110111;
				8'b1000111: c <= 9'b110001;
				8'b1011111: c <= 9'b1100110;
				8'b1110100: c <= 9'b111000011;
				8'b101101: c <= 9'b101110110;
				8'b1010011: c <= 9'b110101111;
				8'b1100001: c <= 9'b101000110;
				8'b110101: c <= 9'b101010101;
				8'b1000100: c <= 9'b101011011;
				8'b1010001: c <= 9'b100011011;
				8'b1010100: c <= 9'b101100110;
				8'b1100110: c <= 9'b10001110;
				8'b101010: c <= 9'b10000010;
				8'b1011110: c <= 9'b101101110;
				8'b1100111: c <= 9'b110011100;
				8'b1011010: c <= 9'b110110101;
				8'b1000010: c <= 9'b100101100;
				8'b111101: c <= 9'b10101111;
				8'b110000: c <= 9'b110100101;
				8'b111110: c <= 9'b101010;
				8'b1100010: c <= 9'b111000100;
				8'b1110000: c <= 9'b110100;
				8'b1101001: c <= 9'b1101010;
				8'b1110011: c <= 9'b111111011;
				8'b1001100: c <= 9'b1011011;
				8'b100001: c <= 9'b100100001;
				8'b1000110: c <= 9'b10110101;
				8'b1110010: c <= 9'b1111111;
				8'b1010000: c <= 9'b10000110;
				8'b1111010: c <= 9'b100011000;
				8'b1010101: c <= 9'b10010001;
				8'b111011: c <= 9'b11100;
				8'b1001101: c <= 9'b101010100;
				8'b111111: c <= 9'b10110011;
				8'b1101110: c <= 9'b100100001;
				8'b1111011: c <= 9'b110110101;
				8'b1001011: c <= 9'b1101;
				8'b1101111: c <= 9'b10111101;
				8'b1101000: c <= 9'b10101001;
				8'b101100: c <= 9'b101001001;
				8'b100100: c <= 9'b1100111;
				8'b1111000: c <= 9'b10000010;
				8'b1000101: c <= 9'b101110001;
				8'b1011001: c <= 9'b110000001;
				8'b110100: c <= 9'b110000000;
				8'b1111001: c <= 9'b11100000;
				8'b1110001: c <= 9'b10100000;
				8'b1001111: c <= 9'b111111111;
				8'b1100101: c <= 9'b111011011;
				8'b1111110: c <= 9'b1111111;
				8'b1111100: c <= 9'b111000000;
				8'b1010110: c <= 9'b100101011;
				8'b110010: c <= 9'b110011101;
				8'b1101101: c <= 9'b11001111;
				8'b100011: c <= 9'b110101;
				8'b1110101: c <= 9'b10011010;
				8'b1111101: c <= 9'b101010001;
				8'b101001: c <= 9'b10111010;
				8'b1010010: c <= 9'b110100111;
				8'b1011000: c <= 9'b1100010;
				8'b101110: c <= 9'b100110010;
				8'b1000001: c <= 9'b110011001;
				default: c <= 9'b0;
			endcase
			9'b100100110 : case(di)
				8'b1000011: c <= 9'b111000101;
				8'b101000: c <= 9'b1100000;
				8'b111010: c <= 9'b11100010;
				8'b110110: c <= 9'b111011001;
				8'b1100100: c <= 9'b101100100;
				8'b1000000: c <= 9'b100101111;
				8'b1110110: c <= 9'b1111111;
				8'b100101: c <= 9'b111101;
				8'b101111: c <= 9'b110101001;
				8'b100110: c <= 9'b100001001;
				8'b1100011: c <= 9'b100010;
				8'b1001000: c <= 9'b10000110;
				8'b111000: c <= 9'b1111101;
				8'b110001: c <= 9'b111000101;
				8'b1010111: c <= 9'b10110101;
				8'b1001110: c <= 9'b1100001;
				8'b1101010: c <= 9'b101001011;
				8'b1001001: c <= 9'b11010101;
				8'b1100000: c <= 9'b1111000;
				8'b110111: c <= 9'b101101000;
				8'b1011101: c <= 9'b111010111;
				8'b1011011: c <= 9'b110;
				8'b111001: c <= 9'b10100100;
				8'b1001010: c <= 9'b110000010;
				8'b110011: c <= 9'b1101;
				8'b1101100: c <= 9'b11111010;
				8'b1110111: c <= 9'b11000011;
				8'b101011: c <= 9'b110010011;
				8'b1101011: c <= 9'b110011100;
				8'b111100: c <= 9'b101100100;
				8'b1000111: c <= 9'b1001110;
				8'b1011111: c <= 9'b10;
				8'b1110100: c <= 9'b1101010;
				8'b101101: c <= 9'b10111101;
				8'b1010011: c <= 9'b101101111;
				8'b1100001: c <= 9'b111111111;
				8'b110101: c <= 9'b111000010;
				8'b1000100: c <= 9'b101000001;
				8'b1010001: c <= 9'b111111001;
				8'b1010100: c <= 9'b10110110;
				8'b1100110: c <= 9'b111111110;
				8'b101010: c <= 9'b111000010;
				8'b1011110: c <= 9'b10001100;
				8'b1100111: c <= 9'b101100100;
				8'b1011010: c <= 9'b11010100;
				8'b1000010: c <= 9'b11010;
				8'b111101: c <= 9'b111111011;
				8'b110000: c <= 9'b110001010;
				8'b111110: c <= 9'b10111;
				8'b1100010: c <= 9'b100000010;
				8'b1110000: c <= 9'b1110111;
				8'b1101001: c <= 9'b100011101;
				8'b1110011: c <= 9'b100010110;
				8'b1001100: c <= 9'b111011010;
				8'b100001: c <= 9'b10111111;
				8'b1000110: c <= 9'b110101111;
				8'b1110010: c <= 9'b110000101;
				8'b1010000: c <= 9'b10100000;
				8'b1111010: c <= 9'b110110111;
				8'b1010101: c <= 9'b1001001;
				8'b111011: c <= 9'b111111;
				8'b1001101: c <= 9'b100000100;
				8'b111111: c <= 9'b11000110;
				8'b1101110: c <= 9'b11;
				8'b1111011: c <= 9'b110111;
				8'b1001011: c <= 9'b100100000;
				8'b1101111: c <= 9'b110001001;
				8'b1101000: c <= 9'b111101001;
				8'b101100: c <= 9'b100010100;
				8'b100100: c <= 9'b111100000;
				8'b1111000: c <= 9'b101110000;
				8'b1000101: c <= 9'b11010111;
				8'b1011001: c <= 9'b110101;
				8'b110100: c <= 9'b110001111;
				8'b1111001: c <= 9'b11011110;
				8'b1110001: c <= 9'b10010111;
				8'b1001111: c <= 9'b1110010;
				8'b1100101: c <= 9'b1000111;
				8'b1111110: c <= 9'b10011001;
				8'b1111100: c <= 9'b101001001;
				8'b1010110: c <= 9'b100000011;
				8'b110010: c <= 9'b101010010;
				8'b1101101: c <= 9'b101110011;
				8'b100011: c <= 9'b100100101;
				8'b1110101: c <= 9'b100100011;
				8'b1111101: c <= 9'b111110011;
				8'b101001: c <= 9'b110100000;
				8'b1010010: c <= 9'b101000111;
				8'b1011000: c <= 9'b101010110;
				8'b101110: c <= 9'b100111000;
				8'b1000001: c <= 9'b110000101;
				default: c <= 9'b0;
			endcase
			9'b10001011 : case(di)
				8'b1000011: c <= 9'b101011010;
				8'b101000: c <= 9'b1101111;
				8'b111010: c <= 9'b110010001;
				8'b110110: c <= 9'b1110000;
				8'b1100100: c <= 9'b11000000;
				8'b1000000: c <= 9'b100110100;
				8'b1110110: c <= 9'b111100111;
				8'b100101: c <= 9'b101110010;
				8'b101111: c <= 9'b101110011;
				8'b100110: c <= 9'b101000;
				8'b1100011: c <= 9'b11000100;
				8'b1001000: c <= 9'b100111000;
				8'b111000: c <= 9'b1111101;
				8'b110001: c <= 9'b111000100;
				8'b1010111: c <= 9'b11110011;
				8'b1001110: c <= 9'b1111101;
				8'b1101010: c <= 9'b100011011;
				8'b1001001: c <= 9'b1010011;
				8'b1100000: c <= 9'b11100;
				8'b110111: c <= 9'b111100011;
				8'b1011101: c <= 9'b101011110;
				8'b1011011: c <= 9'b111001;
				8'b111001: c <= 9'b110111000;
				8'b1001010: c <= 9'b1000101;
				8'b110011: c <= 9'b1011;
				8'b1101100: c <= 9'b100110100;
				8'b1110111: c <= 9'b1111100;
				8'b101011: c <= 9'b1100101;
				8'b1101011: c <= 9'b110010;
				8'b111100: c <= 9'b101100000;
				8'b1000111: c <= 9'b10100;
				8'b1011111: c <= 9'b101101010;
				8'b1110100: c <= 9'b10110011;
				8'b101101: c <= 9'b10100100;
				8'b1010011: c <= 9'b100001010;
				8'b1100001: c <= 9'b100000001;
				8'b110101: c <= 9'b11100111;
				8'b1000100: c <= 9'b11011010;
				8'b1010001: c <= 9'b10010000;
				8'b1010100: c <= 9'b1100011;
				8'b1100110: c <= 9'b10010011;
				8'b101010: c <= 9'b100110011;
				8'b1011110: c <= 9'b10001100;
				8'b1100111: c <= 9'b100011001;
				8'b1011010: c <= 9'b1011110;
				8'b1000010: c <= 9'b110;
				8'b111101: c <= 9'b1100011;
				8'b110000: c <= 9'b10000;
				8'b111110: c <= 9'b110001100;
				8'b1100010: c <= 9'b1010010;
				8'b1110000: c <= 9'b101100111;
				8'b1101001: c <= 9'b100001110;
				8'b1110011: c <= 9'b10000001;
				8'b1001100: c <= 9'b10011100;
				8'b100001: c <= 9'b1000;
				8'b1000110: c <= 9'b111111111;
				8'b1110010: c <= 9'b1011110;
				8'b1010000: c <= 9'b111101111;
				8'b1111010: c <= 9'b1100001;
				8'b1010101: c <= 9'b10011101;
				8'b111011: c <= 9'b110011110;
				8'b1001101: c <= 9'b110010100;
				8'b111111: c <= 9'b101000;
				8'b1101110: c <= 9'b10011111;
				8'b1111011: c <= 9'b100101111;
				8'b1001011: c <= 9'b10100000;
				8'b1101111: c <= 9'b110100010;
				8'b1101000: c <= 9'b10101101;
				8'b101100: c <= 9'b110101010;
				8'b100100: c <= 9'b110101011;
				8'b1111000: c <= 9'b110001001;
				8'b1000101: c <= 9'b111000110;
				8'b1011001: c <= 9'b1001000;
				8'b110100: c <= 9'b111110110;
				8'b1111001: c <= 9'b110011001;
				8'b1110001: c <= 9'b10010001;
				8'b1001111: c <= 9'b100100101;
				8'b1100101: c <= 9'b10011010;
				8'b1111110: c <= 9'b101011011;
				8'b1111100: c <= 9'b111011101;
				8'b1010110: c <= 9'b11110111;
				8'b110010: c <= 9'b10001110;
				8'b1101101: c <= 9'b100100010;
				8'b100011: c <= 9'b1011111;
				8'b1110101: c <= 9'b101000010;
				8'b1111101: c <= 9'b110011100;
				8'b101001: c <= 9'b10111001;
				8'b1010010: c <= 9'b101001111;
				8'b1011000: c <= 9'b101011000;
				8'b101110: c <= 9'b1010010;
				8'b1000001: c <= 9'b10110100;
				default: c <= 9'b0;
			endcase
			9'b10110010 : case(di)
				8'b1000011: c <= 9'b111001111;
				8'b101000: c <= 9'b110011111;
				8'b111010: c <= 9'b101101000;
				8'b110110: c <= 9'b100010111;
				8'b1100100: c <= 9'b11111011;
				8'b1000000: c <= 9'b10001111;
				8'b1110110: c <= 9'b11000000;
				8'b100101: c <= 9'b101100011;
				8'b101111: c <= 9'b1100000;
				8'b100110: c <= 9'b11100010;
				8'b1100011: c <= 9'b111000010;
				8'b1001000: c <= 9'b10101100;
				8'b111000: c <= 9'b10100101;
				8'b110001: c <= 9'b110011000;
				8'b1010111: c <= 9'b11001111;
				8'b1001110: c <= 9'b10001000;
				8'b1101010: c <= 9'b111011011;
				8'b1001001: c <= 9'b101000100;
				8'b1100000: c <= 9'b10000011;
				8'b110111: c <= 9'b101111000;
				8'b1011101: c <= 9'b11111;
				8'b1011011: c <= 9'b111011010;
				8'b111001: c <= 9'b101011101;
				8'b1001010: c <= 9'b110110111;
				8'b110011: c <= 9'b101110;
				8'b1101100: c <= 9'b1110;
				8'b1110111: c <= 9'b11000111;
				8'b101011: c <= 9'b111;
				8'b1101011: c <= 9'b10010100;
				8'b111100: c <= 9'b1111101;
				8'b1000111: c <= 9'b11101111;
				8'b1011111: c <= 9'b10011;
				8'b1110100: c <= 9'b1101000;
				8'b101101: c <= 9'b111011;
				8'b1010011: c <= 9'b1;
				8'b1100001: c <= 9'b11110;
				8'b110101: c <= 9'b111100000;
				8'b1000100: c <= 9'b1111010;
				8'b1010001: c <= 9'b100110000;
				8'b1010100: c <= 9'b10010001;
				8'b1100110: c <= 9'b111010110;
				8'b101010: c <= 9'b111101;
				8'b1011110: c <= 9'b10010011;
				8'b1100111: c <= 9'b11001010;
				8'b1011010: c <= 9'b111000110;
				8'b1000010: c <= 9'b101100011;
				8'b111101: c <= 9'b1110010;
				8'b110000: c <= 9'b11000110;
				8'b111110: c <= 9'b10111111;
				8'b1100010: c <= 9'b100001110;
				8'b1110000: c <= 9'b10011;
				8'b1101001: c <= 9'b110010;
				8'b1110011: c <= 9'b111001010;
				8'b1001100: c <= 9'b1100111;
				8'b100001: c <= 9'b100000011;
				8'b1000110: c <= 9'b101111000;
				8'b1110010: c <= 9'b11011;
				8'b1010000: c <= 9'b101010;
				8'b1111010: c <= 9'b11011;
				8'b1010101: c <= 9'b10101011;
				8'b111011: c <= 9'b101010010;
				8'b1001101: c <= 9'b110100;
				8'b111111: c <= 9'b101101010;
				8'b1101110: c <= 9'b10110010;
				8'b1111011: c <= 9'b100111111;
				8'b1001011: c <= 9'b100111001;
				8'b1101111: c <= 9'b110010;
				8'b1101000: c <= 9'b110110011;
				8'b101100: c <= 9'b10000010;
				8'b100100: c <= 9'b111011001;
				8'b1111000: c <= 9'b10101110;
				8'b1000101: c <= 9'b111001001;
				8'b1011001: c <= 9'b110000000;
				8'b110100: c <= 9'b110001100;
				8'b1111001: c <= 9'b1000001;
				8'b1110001: c <= 9'b111011;
				8'b1001111: c <= 9'b110011;
				8'b1100101: c <= 9'b11110110;
				8'b1111110: c <= 9'b100000100;
				8'b1111100: c <= 9'b1101;
				8'b1010110: c <= 9'b1010000;
				8'b110010: c <= 9'b100100101;
				8'b1101101: c <= 9'b11110101;
				8'b100011: c <= 9'b1010001;
				8'b1110101: c <= 9'b1101100;
				8'b1111101: c <= 9'b1001000;
				8'b101001: c <= 9'b100010001;
				8'b1010010: c <= 9'b1111;
				8'b1011000: c <= 9'b10110011;
				8'b101110: c <= 9'b10101101;
				8'b1000001: c <= 9'b100001111;
				default: c <= 9'b0;
			endcase
			9'b11101001 : case(di)
				8'b1000011: c <= 9'b1010010;
				8'b101000: c <= 9'b100100001;
				8'b111010: c <= 9'b110001;
				8'b110110: c <= 9'b101010100;
				8'b1100100: c <= 9'b101;
				8'b1000000: c <= 9'b110000111;
				8'b1110110: c <= 9'b101101111;
				8'b100101: c <= 9'b10011001;
				8'b101111: c <= 9'b101001;
				8'b100110: c <= 9'b110000000;
				8'b1100011: c <= 9'b1011100;
				8'b1001000: c <= 9'b100110000;
				8'b111000: c <= 9'b101100010;
				8'b110001: c <= 9'b11011;
				8'b1010111: c <= 9'b111111000;
				8'b1001110: c <= 9'b111;
				8'b1101010: c <= 9'b111000110;
				8'b1001001: c <= 9'b1000010;
				8'b1100000: c <= 9'b110000101;
				8'b110111: c <= 9'b110010010;
				8'b1011101: c <= 9'b11110;
				8'b1011011: c <= 9'b10111110;
				8'b111001: c <= 9'b10100010;
				8'b1001010: c <= 9'b101101100;
				8'b110011: c <= 9'b1010111;
				8'b1101100: c <= 9'b1000000;
				8'b1110111: c <= 9'b10001011;
				8'b101011: c <= 9'b110001101;
				8'b1101011: c <= 9'b111111011;
				8'b111100: c <= 9'b1111000;
				8'b1000111: c <= 9'b101110101;
				8'b1011111: c <= 9'b11111011;
				8'b1110100: c <= 9'b111100101;
				8'b101101: c <= 9'b100000110;
				8'b1010011: c <= 9'b111111111;
				8'b1100001: c <= 9'b1101;
				8'b110101: c <= 9'b11010111;
				8'b1000100: c <= 9'b1100001;
				8'b1010001: c <= 9'b11000010;
				8'b1010100: c <= 9'b10000000;
				8'b1100110: c <= 9'b101101001;
				8'b101010: c <= 9'b11100100;
				8'b1011110: c <= 9'b11100000;
				8'b1100111: c <= 9'b100001;
				8'b1011010: c <= 9'b110100100;
				8'b1000010: c <= 9'b1111000;
				8'b111101: c <= 9'b11010001;
				8'b110000: c <= 9'b11000000;
				8'b111110: c <= 9'b110101001;
				8'b1100010: c <= 9'b10011101;
				8'b1110000: c <= 9'b101101101;
				8'b1101001: c <= 9'b101000111;
				8'b1110011: c <= 9'b100011000;
				8'b1001100: c <= 9'b111101100;
				8'b100001: c <= 9'b111111000;
				8'b1000110: c <= 9'b11110011;
				8'b1110010: c <= 9'b111011100;
				8'b1010000: c <= 9'b100000111;
				8'b1111010: c <= 9'b10101;
				8'b1010101: c <= 9'b100100000;
				8'b111011: c <= 9'b10101011;
				8'b1001101: c <= 9'b1111110;
				8'b111111: c <= 9'b101010000;
				8'b1101110: c <= 9'b100101110;
				8'b1111011: c <= 9'b101011101;
				8'b1001011: c <= 9'b101111110;
				8'b1101111: c <= 9'b101100001;
				8'b1101000: c <= 9'b1100101;
				8'b101100: c <= 9'b1100011;
				8'b100100: c <= 9'b111100110;
				8'b1111000: c <= 9'b100001;
				8'b1000101: c <= 9'b110101010;
				8'b1011001: c <= 9'b1101100;
				8'b110100: c <= 9'b11010101;
				8'b1111001: c <= 9'b110010100;
				8'b1110001: c <= 9'b11111011;
				8'b1001111: c <= 9'b110110101;
				8'b1100101: c <= 9'b10000101;
				8'b1111110: c <= 9'b101010101;
				8'b1111100: c <= 9'b1100001;
				8'b1010110: c <= 9'b100000001;
				8'b110010: c <= 9'b110100110;
				8'b1101101: c <= 9'b1010011;
				8'b100011: c <= 9'b1110000;
				8'b1110101: c <= 9'b100100101;
				8'b1111101: c <= 9'b110101011;
				8'b101001: c <= 9'b10011011;
				8'b1010010: c <= 9'b101100001;
				8'b1011000: c <= 9'b10101000;
				8'b101110: c <= 9'b11001;
				8'b1000001: c <= 9'b101001000;
				default: c <= 9'b0;
			endcase
			9'b110110101 : case(di)
				8'b1000011: c <= 9'b100010;
				8'b101000: c <= 9'b101100101;
				8'b111010: c <= 9'b1000;
				8'b110110: c <= 9'b111011111;
				8'b1100100: c <= 9'b10000010;
				8'b1000000: c <= 9'b100100111;
				8'b1110110: c <= 9'b1101111;
				8'b100101: c <= 9'b11000111;
				8'b101111: c <= 9'b101000011;
				8'b100110: c <= 9'b10100101;
				8'b1100011: c <= 9'b10001101;
				8'b1001000: c <= 9'b110100010;
				8'b111000: c <= 9'b11110000;
				8'b110001: c <= 9'b1000110;
				8'b1010111: c <= 9'b101000110;
				8'b1001110: c <= 9'b110011100;
				8'b1101010: c <= 9'b11001100;
				8'b1001001: c <= 9'b1010101;
				8'b1100000: c <= 9'b110011100;
				8'b110111: c <= 9'b10;
				8'b1011101: c <= 9'b10;
				8'b1011011: c <= 9'b101101;
				8'b111001: c <= 9'b100110100;
				8'b1001010: c <= 9'b110100001;
				8'b110011: c <= 9'b10101;
				8'b1101100: c <= 9'b11010001;
				8'b1110111: c <= 9'b100111111;
				8'b101011: c <= 9'b10101101;
				8'b1101011: c <= 9'b110;
				8'b111100: c <= 9'b110011101;
				8'b1000111: c <= 9'b110010001;
				8'b1011111: c <= 9'b11111001;
				8'b1110100: c <= 9'b11110010;
				8'b101101: c <= 9'b10111011;
				8'b1010011: c <= 9'b101101100;
				8'b1100001: c <= 9'b11101;
				8'b110101: c <= 9'b101000;
				8'b1000100: c <= 9'b10010000;
				8'b1010001: c <= 9'b111111011;
				8'b1010100: c <= 9'b101101011;
				8'b1100110: c <= 9'b111110101;
				8'b101010: c <= 9'b10110001;
				8'b1011110: c <= 9'b11000;
				8'b1100111: c <= 9'b11000;
				8'b1011010: c <= 9'b100000101;
				8'b1000010: c <= 9'b110001111;
				8'b111101: c <= 9'b111001011;
				8'b110000: c <= 9'b100111100;
				8'b111110: c <= 9'b1010010;
				8'b1100010: c <= 9'b110110010;
				8'b1110000: c <= 9'b10111110;
				8'b1101001: c <= 9'b101101011;
				8'b1110011: c <= 9'b101110011;
				8'b1001100: c <= 9'b110111001;
				8'b100001: c <= 9'b111110011;
				8'b1000110: c <= 9'b100011001;
				8'b1110010: c <= 9'b100111000;
				8'b1010000: c <= 9'b1010010;
				8'b1111010: c <= 9'b100010;
				8'b1010101: c <= 9'b10001000;
				8'b111011: c <= 9'b111101101;
				8'b1001101: c <= 9'b111100110;
				8'b111111: c <= 9'b1010111;
				8'b1101110: c <= 9'b11000000;
				8'b1111011: c <= 9'b111000010;
				8'b1001011: c <= 9'b11010100;
				8'b1101111: c <= 9'b100010110;
				8'b1101000: c <= 9'b10011;
				8'b101100: c <= 9'b100001101;
				8'b100100: c <= 9'b111000;
				8'b1111000: c <= 9'b110010010;
				8'b1000101: c <= 9'b110001001;
				8'b1011001: c <= 9'b11110010;
				8'b110100: c <= 9'b1110011;
				8'b1111001: c <= 9'b111000100;
				8'b1110001: c <= 9'b101110110;
				8'b1001111: c <= 9'b101111111;
				8'b1100101: c <= 9'b100011001;
				8'b1111110: c <= 9'b10101110;
				8'b1111100: c <= 9'b10010011;
				8'b1010110: c <= 9'b10100;
				8'b110010: c <= 9'b101100101;
				8'b1101101: c <= 9'b1000;
				8'b100011: c <= 9'b101101011;
				8'b1110101: c <= 9'b111001010;
				8'b1111101: c <= 9'b101110001;
				8'b101001: c <= 9'b111010000;
				8'b1010010: c <= 9'b111010;
				8'b1011000: c <= 9'b111001101;
				8'b101110: c <= 9'b1111111;
				8'b1000001: c <= 9'b11101100;
				default: c <= 9'b0;
			endcase
			9'b100000111 : case(di)
				8'b1000011: c <= 9'b10101100;
				8'b101000: c <= 9'b101100010;
				8'b111010: c <= 9'b101001010;
				8'b110110: c <= 9'b1010010;
				8'b1100100: c <= 9'b100111010;
				8'b1000000: c <= 9'b111101110;
				8'b1110110: c <= 9'b110000000;
				8'b100101: c <= 9'b111001101;
				8'b101111: c <= 9'b10011010;
				8'b100110: c <= 9'b11001010;
				8'b1100011: c <= 9'b110011;
				8'b1001000: c <= 9'b10000010;
				8'b111000: c <= 9'b100001010;
				8'b110001: c <= 9'b100001011;
				8'b1010111: c <= 9'b11100011;
				8'b1001110: c <= 9'b110101;
				8'b1101010: c <= 9'b110101110;
				8'b1001001: c <= 9'b110011101;
				8'b1100000: c <= 9'b11110110;
				8'b110111: c <= 9'b110111001;
				8'b1011101: c <= 9'b101101;
				8'b1011011: c <= 9'b101001010;
				8'b111001: c <= 9'b111100101;
				8'b1001010: c <= 9'b11100000;
				8'b110011: c <= 9'b10110011;
				8'b1101100: c <= 9'b11100111;
				8'b1110111: c <= 9'b100111000;
				8'b101011: c <= 9'b111110101;
				8'b1101011: c <= 9'b100010000;
				8'b111100: c <= 9'b101100;
				8'b1000111: c <= 9'b101001010;
				8'b1011111: c <= 9'b10011010;
				8'b1110100: c <= 9'b110111;
				8'b101101: c <= 9'b10000011;
				8'b1010011: c <= 9'b100111010;
				8'b1100001: c <= 9'b100011001;
				8'b110101: c <= 9'b110111011;
				8'b1000100: c <= 9'b111001;
				8'b1010001: c <= 9'b111001011;
				8'b1010100: c <= 9'b110101110;
				8'b1100110: c <= 9'b101011110;
				8'b101010: c <= 9'b1010111;
				8'b1011110: c <= 9'b101101010;
				8'b1100111: c <= 9'b101100111;
				8'b1011010: c <= 9'b11011000;
				8'b1000010: c <= 9'b11100010;
				8'b111101: c <= 9'b101011;
				8'b110000: c <= 9'b11011110;
				8'b111110: c <= 9'b11011001;
				8'b1100010: c <= 9'b110001000;
				8'b1110000: c <= 9'b100000111;
				8'b1101001: c <= 9'b110111001;
				8'b1110011: c <= 9'b110010111;
				8'b1001100: c <= 9'b111010;
				8'b100001: c <= 9'b101001;
				8'b1000110: c <= 9'b100010110;
				8'b1110010: c <= 9'b100011000;
				8'b1010000: c <= 9'b1101010;
				8'b1111010: c <= 9'b111000;
				8'b1010101: c <= 9'b110001;
				8'b111011: c <= 9'b100001100;
				8'b1001101: c <= 9'b1110000;
				8'b111111: c <= 9'b111101;
				8'b1101110: c <= 9'b10001001;
				8'b1111011: c <= 9'b100110111;
				8'b1001011: c <= 9'b11011011;
				8'b1101111: c <= 9'b110000001;
				8'b1101000: c <= 9'b110000011;
				8'b101100: c <= 9'b110101001;
				8'b100100: c <= 9'b100110100;
				8'b1111000: c <= 9'b100001010;
				8'b1000101: c <= 9'b100010100;
				8'b1011001: c <= 9'b10011010;
				8'b110100: c <= 9'b10001111;
				8'b1111001: c <= 9'b10111100;
				8'b1110001: c <= 9'b111000000;
				8'b1001111: c <= 9'b100000000;
				8'b1100101: c <= 9'b100010100;
				8'b1111110: c <= 9'b101110101;
				8'b1111100: c <= 9'b110001001;
				8'b1010110: c <= 9'b1000;
				8'b110010: c <= 9'b100000101;
				8'b1101101: c <= 9'b11100100;
				8'b100011: c <= 9'b101001010;
				8'b1110101: c <= 9'b10000101;
				8'b1111101: c <= 9'b111000100;
				8'b101001: c <= 9'b1010111;
				8'b1010010: c <= 9'b101000;
				8'b1011000: c <= 9'b1111101;
				8'b101110: c <= 9'b11110001;
				8'b1000001: c <= 9'b110011001;
				default: c <= 9'b0;
			endcase
			9'b110010101 : case(di)
				8'b1000011: c <= 9'b110100000;
				8'b101000: c <= 9'b111001101;
				8'b111010: c <= 9'b111001100;
				8'b110110: c <= 9'b100000111;
				8'b1100100: c <= 9'b101000110;
				8'b1000000: c <= 9'b110000011;
				8'b1110110: c <= 9'b110110111;
				8'b100101: c <= 9'b100001101;
				8'b101111: c <= 9'b101010000;
				8'b100110: c <= 9'b110000110;
				8'b1100011: c <= 9'b100111000;
				8'b1001000: c <= 9'b10000010;
				8'b111000: c <= 9'b110001101;
				8'b110001: c <= 9'b101101010;
				8'b1010111: c <= 9'b10111101;
				8'b1001110: c <= 9'b111011110;
				8'b1101010: c <= 9'b110001111;
				8'b1001001: c <= 9'b100111101;
				8'b1100000: c <= 9'b10000110;
				8'b110111: c <= 9'b101101001;
				8'b1011101: c <= 9'b11100101;
				8'b1011011: c <= 9'b10101110;
				8'b111001: c <= 9'b100;
				8'b1001010: c <= 9'b110111100;
				8'b110011: c <= 9'b111100111;
				8'b1101100: c <= 9'b100010010;
				8'b1110111: c <= 9'b110110011;
				8'b101011: c <= 9'b101010011;
				8'b1101011: c <= 9'b111001011;
				8'b111100: c <= 9'b100111000;
				8'b1000111: c <= 9'b10110001;
				8'b1011111: c <= 9'b11110101;
				8'b1110100: c <= 9'b1001000;
				8'b101101: c <= 9'b101101100;
				8'b1010011: c <= 9'b110001100;
				8'b1100001: c <= 9'b100101011;
				8'b110101: c <= 9'b110000111;
				8'b1000100: c <= 9'b101001;
				8'b1010001: c <= 9'b10101010;
				8'b1010100: c <= 9'b11111010;
				8'b1100110: c <= 9'b110011;
				8'b101010: c <= 9'b10010001;
				8'b1011110: c <= 9'b110001111;
				8'b1100111: c <= 9'b111111001;
				8'b1011010: c <= 9'b100010000;
				8'b1000010: c <= 9'b101000001;
				8'b111101: c <= 9'b10000000;
				8'b110000: c <= 9'b10111110;
				8'b111110: c <= 9'b100101010;
				8'b1100010: c <= 9'b110000011;
				8'b1110000: c <= 9'b101001111;
				8'b1101001: c <= 9'b101100011;
				8'b1110011: c <= 9'b100111010;
				8'b1001100: c <= 9'b111000101;
				8'b100001: c <= 9'b10001101;
				8'b1000110: c <= 9'b1110100;
				8'b1110010: c <= 9'b1001111;
				8'b1010000: c <= 9'b10110110;
				8'b1111010: c <= 9'b111010110;
				8'b1010101: c <= 9'b101110111;
				8'b111011: c <= 9'b100110101;
				8'b1001101: c <= 9'b101010011;
				8'b111111: c <= 9'b101000111;
				8'b1101110: c <= 9'b100001101;
				8'b1111011: c <= 9'b10111;
				8'b1001011: c <= 9'b100111000;
				8'b1101111: c <= 9'b10001100;
				8'b1101000: c <= 9'b101001110;
				8'b101100: c <= 9'b11000100;
				8'b100100: c <= 9'b111111011;
				8'b1111000: c <= 9'b111010010;
				8'b1000101: c <= 9'b101101111;
				8'b1011001: c <= 9'b110010011;
				8'b110100: c <= 9'b10010110;
				8'b1111001: c <= 9'b1100011;
				8'b1110001: c <= 9'b100101101;
				8'b1001111: c <= 9'b111100;
				8'b1100101: c <= 9'b110001010;
				8'b1111110: c <= 9'b10011010;
				8'b1111100: c <= 9'b111111000;
				8'b1010110: c <= 9'b101000;
				8'b110010: c <= 9'b101101111;
				8'b1101101: c <= 9'b10011001;
				8'b100011: c <= 9'b11100000;
				8'b1110101: c <= 9'b10100100;
				8'b1111101: c <= 9'b10111000;
				8'b101001: c <= 9'b101011;
				8'b1010010: c <= 9'b10100011;
				8'b1011000: c <= 9'b10101111;
				8'b101110: c <= 9'b11110;
				8'b1000001: c <= 9'b10101000;
				default: c <= 9'b0;
			endcase
			9'b100010101 : case(di)
				8'b1000011: c <= 9'b101110101;
				8'b101000: c <= 9'b10001001;
				8'b111010: c <= 9'b110101001;
				8'b110110: c <= 9'b101001000;
				8'b1100100: c <= 9'b10111001;
				8'b1000000: c <= 9'b111101000;
				8'b1110110: c <= 9'b110110111;
				8'b100101: c <= 9'b110010110;
				8'b101111: c <= 9'b1011110;
				8'b100110: c <= 9'b10011010;
				8'b1100011: c <= 9'b101011111;
				8'b1001000: c <= 9'b11000111;
				8'b111000: c <= 9'b100001111;
				8'b110001: c <= 9'b111100111;
				8'b1010111: c <= 9'b110100101;
				8'b1001110: c <= 9'b1101010;
				8'b1101010: c <= 9'b1100;
				8'b1001001: c <= 9'b1110001;
				8'b1100000: c <= 9'b10100100;
				8'b110111: c <= 9'b1111101;
				8'b1011101: c <= 9'b110;
				8'b1011011: c <= 9'b11011;
				8'b111001: c <= 9'b110111010;
				8'b1001010: c <= 9'b111010000;
				8'b110011: c <= 9'b100111101;
				8'b1101100: c <= 9'b110101101;
				8'b1110111: c <= 9'b101100;
				8'b101011: c <= 9'b11111000;
				8'b1101011: c <= 9'b110111111;
				8'b111100: c <= 9'b110110011;
				8'b1000111: c <= 9'b10101100;
				8'b1011111: c <= 9'b10101010;
				8'b1110100: c <= 9'b10000001;
				8'b101101: c <= 9'b100010110;
				8'b1010011: c <= 9'b110010001;
				8'b1100001: c <= 9'b1011111;
				8'b110101: c <= 9'b10101;
				8'b1000100: c <= 9'b110100011;
				8'b1010001: c <= 9'b11011100;
				8'b1010100: c <= 9'b10000001;
				8'b1100110: c <= 9'b100010110;
				8'b101010: c <= 9'b101111010;
				8'b1011110: c <= 9'b11000;
				8'b1100111: c <= 9'b110111011;
				8'b1011010: c <= 9'b100101010;
				8'b1000010: c <= 9'b111101110;
				8'b111101: c <= 9'b100110010;
				8'b110000: c <= 9'b111100100;
				8'b111110: c <= 9'b10100010;
				8'b1100010: c <= 9'b110111100;
				8'b1110000: c <= 9'b10101110;
				8'b1101001: c <= 9'b110000001;
				8'b1110011: c <= 9'b110101111;
				8'b1001100: c <= 9'b101011000;
				8'b100001: c <= 9'b1100110;
				8'b1000110: c <= 9'b110100100;
				8'b1110010: c <= 9'b111001010;
				8'b1010000: c <= 9'b110011;
				8'b1111010: c <= 9'b1011111;
				8'b1010101: c <= 9'b110110100;
				8'b111011: c <= 9'b100101;
				8'b1001101: c <= 9'b10011100;
				8'b111111: c <= 9'b100110101;
				8'b1101110: c <= 9'b1000111;
				8'b1111011: c <= 9'b11000000;
				8'b1001011: c <= 9'b100001101;
				8'b1101111: c <= 9'b100000000;
				8'b1101000: c <= 9'b11100011;
				8'b101100: c <= 9'b100111001;
				8'b100100: c <= 9'b100010000;
				8'b1111000: c <= 9'b101000;
				8'b1000101: c <= 9'b100111011;
				8'b1011001: c <= 9'b10001101;
				8'b110100: c <= 9'b111010001;
				8'b1111001: c <= 9'b100110111;
				8'b1110001: c <= 9'b100110000;
				8'b1001111: c <= 9'b100110100;
				8'b1100101: c <= 9'b101010;
				8'b1111110: c <= 9'b100100001;
				8'b1111100: c <= 9'b1100111;
				8'b1010110: c <= 9'b110111011;
				8'b110010: c <= 9'b111010000;
				8'b1101101: c <= 9'b1000110;
				8'b100011: c <= 9'b10101110;
				8'b1110101: c <= 9'b101101111;
				8'b1111101: c <= 9'b100101010;
				8'b101001: c <= 9'b100000010;
				8'b1010010: c <= 9'b10101100;
				8'b1011000: c <= 9'b111101010;
				8'b101110: c <= 9'b111011;
				8'b1000001: c <= 9'b101000;
				default: c <= 9'b0;
			endcase
			9'b111101110 : case(di)
				8'b1000011: c <= 9'b10100101;
				8'b101000: c <= 9'b100101000;
				8'b111010: c <= 9'b11010100;
				8'b110110: c <= 9'b110111111;
				8'b1100100: c <= 9'b1001001;
				8'b1000000: c <= 9'b100101000;
				8'b1110110: c <= 9'b1100011;
				8'b100101: c <= 9'b110101011;
				8'b101111: c <= 9'b110000111;
				8'b100110: c <= 9'b110111000;
				8'b1100011: c <= 9'b111100010;
				8'b1001000: c <= 9'b111100111;
				8'b111000: c <= 9'b101110111;
				8'b110001: c <= 9'b101011010;
				8'b1010111: c <= 9'b110101011;
				8'b1001110: c <= 9'b110100001;
				8'b1101010: c <= 9'b1100010;
				8'b1001001: c <= 9'b11001;
				8'b1100000: c <= 9'b110101100;
				8'b110111: c <= 9'b11010;
				8'b1011101: c <= 9'b1110001;
				8'b1011011: c <= 9'b1001101;
				8'b111001: c <= 9'b10011111;
				8'b1001010: c <= 9'b111110000;
				8'b110011: c <= 9'b1011100;
				8'b1101100: c <= 9'b11011100;
				8'b1110111: c <= 9'b101001000;
				8'b101011: c <= 9'b110010011;
				8'b1101011: c <= 9'b100111111;
				8'b111100: c <= 9'b10100110;
				8'b1000111: c <= 9'b11101100;
				8'b1011111: c <= 9'b101110000;
				8'b1110100: c <= 9'b11011100;
				8'b101101: c <= 9'b11000110;
				8'b1010011: c <= 9'b10010001;
				8'b1100001: c <= 9'b101000110;
				8'b110101: c <= 9'b101101111;
				8'b1000100: c <= 9'b1110;
				8'b1010001: c <= 9'b1001001;
				8'b1010100: c <= 9'b111100000;
				8'b1100110: c <= 9'b11001101;
				8'b101010: c <= 9'b100011101;
				8'b1011110: c <= 9'b100110100;
				8'b1100111: c <= 9'b100001100;
				8'b1011010: c <= 9'b101000110;
				8'b1000010: c <= 9'b1010110;
				8'b111101: c <= 9'b100011000;
				8'b110000: c <= 9'b100011011;
				8'b111110: c <= 9'b10110;
				8'b1100010: c <= 9'b11110101;
				8'b1110000: c <= 9'b100110101;
				8'b1101001: c <= 9'b10101101;
				8'b1110011: c <= 9'b110101011;
				8'b1001100: c <= 9'b101111010;
				8'b100001: c <= 9'b10011101;
				8'b1000110: c <= 9'b100010110;
				8'b1110010: c <= 9'b110111110;
				8'b1010000: c <= 9'b1001110;
				8'b1111010: c <= 9'b10110101;
				8'b1010101: c <= 9'b1000100;
				8'b111011: c <= 9'b11110;
				8'b1001101: c <= 9'b111001010;
				8'b111111: c <= 9'b101101110;
				8'b1101110: c <= 9'b100001001;
				8'b1111011: c <= 9'b10100000;
				8'b1001011: c <= 9'b1101110;
				8'b1101111: c <= 9'b101010;
				8'b1101000: c <= 9'b1010110;
				8'b101100: c <= 9'b10000111;
				8'b100100: c <= 9'b111000101;
				8'b1111000: c <= 9'b101001;
				8'b1000101: c <= 9'b1110010;
				8'b1011001: c <= 9'b100110;
				8'b110100: c <= 9'b100101010;
				8'b1111001: c <= 9'b10110111;
				8'b1110001: c <= 9'b101011000;
				8'b1001111: c <= 9'b1100011;
				8'b1100101: c <= 9'b1100011;
				8'b1111110: c <= 9'b110111100;
				8'b1111100: c <= 9'b1111100;
				8'b1010110: c <= 9'b10001011;
				8'b110010: c <= 9'b111001010;
				8'b1101101: c <= 9'b1101010;
				8'b100011: c <= 9'b110000010;
				8'b1110101: c <= 9'b11010010;
				8'b1111101: c <= 9'b110100110;
				8'b101001: c <= 9'b101001011;
				8'b1010010: c <= 9'b11100001;
				8'b1011000: c <= 9'b100001110;
				8'b101110: c <= 9'b10000000;
				8'b1000001: c <= 9'b11101001;
				default: c <= 9'b0;
			endcase
			9'b100001011 : case(di)
				8'b1000011: c <= 9'b100111011;
				8'b101000: c <= 9'b10110100;
				8'b111010: c <= 9'b111010010;
				8'b110110: c <= 9'b110000;
				8'b1100100: c <= 9'b1001110;
				8'b1000000: c <= 9'b10100000;
				8'b1110110: c <= 9'b1101000;
				8'b100101: c <= 9'b1001100;
				8'b101111: c <= 9'b10010101;
				8'b100110: c <= 9'b101000111;
				8'b1100011: c <= 9'b110110000;
				8'b1001000: c <= 9'b10001100;
				8'b111000: c <= 9'b101000110;
				8'b110001: c <= 9'b1110011;
				8'b1010111: c <= 9'b101111111;
				8'b1001110: c <= 9'b1110;
				8'b1101010: c <= 9'b111111101;
				8'b1001001: c <= 9'b101111110;
				8'b1100000: c <= 9'b100111101;
				8'b110111: c <= 9'b110110110;
				8'b1011101: c <= 9'b101101;
				8'b1011011: c <= 9'b101111000;
				8'b111001: c <= 9'b101011011;
				8'b1001010: c <= 9'b10010011;
				8'b110011: c <= 9'b1011100;
				8'b1101100: c <= 9'b10110101;
				8'b1110111: c <= 9'b101100111;
				8'b101011: c <= 9'b110010001;
				8'b1101011: c <= 9'b11110001;
				8'b111100: c <= 9'b101010100;
				8'b1000111: c <= 9'b1111010;
				8'b1011111: c <= 9'b100000011;
				8'b1110100: c <= 9'b100010101;
				8'b101101: c <= 9'b110110011;
				8'b1010011: c <= 9'b111111001;
				8'b1100001: c <= 9'b1000111;
				8'b110101: c <= 9'b101011000;
				8'b1000100: c <= 9'b110111;
				8'b1010001: c <= 9'b110011011;
				8'b1010100: c <= 9'b1100;
				8'b1100110: c <= 9'b101011001;
				8'b101010: c <= 9'b11010100;
				8'b1011110: c <= 9'b111001011;
				8'b1100111: c <= 9'b110011110;
				8'b1011010: c <= 9'b1111101;
				8'b1000010: c <= 9'b111110001;
				8'b111101: c <= 9'b111010100;
				8'b110000: c <= 9'b11111100;
				8'b111110: c <= 9'b101110010;
				8'b1100010: c <= 9'b11001000;
				8'b1110000: c <= 9'b10;
				8'b1101001: c <= 9'b101100100;
				8'b1110011: c <= 9'b100000001;
				8'b1001100: c <= 9'b111111101;
				8'b100001: c <= 9'b110001111;
				8'b1000110: c <= 9'b1100001;
				8'b1110010: c <= 9'b100011111;
				8'b1010000: c <= 9'b100101111;
				8'b1111010: c <= 9'b110000110;
				8'b1010101: c <= 9'b1010001;
				8'b111011: c <= 9'b101010001;
				8'b1001101: c <= 9'b1011100;
				8'b111111: c <= 9'b100100110;
				8'b1101110: c <= 9'b10001010;
				8'b1111011: c <= 9'b110011000;
				8'b1001011: c <= 9'b110100101;
				8'b1101111: c <= 9'b111011001;
				8'b1101000: c <= 9'b111100110;
				8'b101100: c <= 9'b110001100;
				8'b100100: c <= 9'b100011000;
				8'b1111000: c <= 9'b10011101;
				8'b1000101: c <= 9'b111010;
				8'b1011001: c <= 9'b101001;
				8'b110100: c <= 9'b110110;
				8'b1111001: c <= 9'b101001011;
				8'b1110001: c <= 9'b10011;
				8'b1001111: c <= 9'b11001100;
				8'b1100101: c <= 9'b1100101;
				8'b1111110: c <= 9'b100110011;
				8'b1111100: c <= 9'b11000000;
				8'b1010110: c <= 9'b10011000;
				8'b110010: c <= 9'b110000000;
				8'b1101101: c <= 9'b10;
				8'b100011: c <= 9'b100011100;
				8'b1110101: c <= 9'b100111001;
				8'b1111101: c <= 9'b11010011;
				8'b101001: c <= 9'b1;
				8'b1010010: c <= 9'b110010101;
				8'b1011000: c <= 9'b11011110;
				8'b101110: c <= 9'b100110101;
				8'b1000001: c <= 9'b10110010;
				default: c <= 9'b0;
			endcase
			9'b100110100 : case(di)
				8'b1000011: c <= 9'b101000101;
				8'b101000: c <= 9'b111011011;
				8'b111010: c <= 9'b1000111;
				8'b110110: c <= 9'b10010101;
				8'b1100100: c <= 9'b111000011;
				8'b1000000: c <= 9'b11100;
				8'b1110110: c <= 9'b111010010;
				8'b100101: c <= 9'b11000111;
				8'b101111: c <= 9'b10001001;
				8'b100110: c <= 9'b101010011;
				8'b1100011: c <= 9'b100101;
				8'b1001000: c <= 9'b10000001;
				8'b111000: c <= 9'b1001001;
				8'b110001: c <= 9'b111100001;
				8'b1010111: c <= 9'b1010000;
				8'b1001110: c <= 9'b11100111;
				8'b1101010: c <= 9'b100101100;
				8'b1001001: c <= 9'b101110;
				8'b1100000: c <= 9'b110010100;
				8'b110111: c <= 9'b111011;
				8'b1011101: c <= 9'b11011010;
				8'b1011011: c <= 9'b10110010;
				8'b111001: c <= 9'b101001110;
				8'b1001010: c <= 9'b110100010;
				8'b110011: c <= 9'b11010;
				8'b1101100: c <= 9'b101110110;
				8'b1110111: c <= 9'b100101000;
				8'b101011: c <= 9'b1110;
				8'b1101011: c <= 9'b111111001;
				8'b111100: c <= 9'b10010;
				8'b1000111: c <= 9'b100101100;
				8'b1011111: c <= 9'b111010110;
				8'b1110100: c <= 9'b10001000;
				8'b101101: c <= 9'b110011;
				8'b1010011: c <= 9'b10100000;
				8'b1100001: c <= 9'b100101100;
				8'b110101: c <= 9'b101011000;
				8'b1000100: c <= 9'b1011;
				8'b1010001: c <= 9'b10001011;
				8'b1010100: c <= 9'b100010110;
				8'b1100110: c <= 9'b10010111;
				8'b101010: c <= 9'b100100101;
				8'b1011110: c <= 9'b110101;
				8'b1100111: c <= 9'b111111;
				8'b1011010: c <= 9'b10111000;
				8'b1000010: c <= 9'b101100001;
				8'b111101: c <= 9'b101000111;
				8'b110000: c <= 9'b100001011;
				8'b111110: c <= 9'b11101101;
				8'b1100010: c <= 9'b101001001;
				8'b1110000: c <= 9'b100000010;
				8'b1101001: c <= 9'b1101000;
				8'b1110011: c <= 9'b101101011;
				8'b1001100: c <= 9'b101100;
				8'b100001: c <= 9'b101000101;
				8'b1000110: c <= 9'b111111111;
				8'b1110010: c <= 9'b10010011;
				8'b1010000: c <= 9'b10100011;
				8'b1111010: c <= 9'b11110111;
				8'b1010101: c <= 9'b1011001;
				8'b111011: c <= 9'b100100111;
				8'b1001101: c <= 9'b11101001;
				8'b111111: c <= 9'b111111101;
				8'b1101110: c <= 9'b11101100;
				8'b1111011: c <= 9'b1111101;
				8'b1001011: c <= 9'b101011110;
				8'b1101111: c <= 9'b11110000;
				8'b1101000: c <= 9'b1101;
				8'b101100: c <= 9'b1111010;
				8'b100100: c <= 9'b11001111;
				8'b1111000: c <= 9'b100011011;
				8'b1000101: c <= 9'b10100010;
				8'b1011001: c <= 9'b110010100;
				8'b110100: c <= 9'b10010000;
				8'b1111001: c <= 9'b10011000;
				8'b1110001: c <= 9'b11000110;
				8'b1001111: c <= 9'b110110111;
				8'b1100101: c <= 9'b110000000;
				8'b1111110: c <= 9'b101100010;
				8'b1111100: c <= 9'b11011000;
				8'b1010110: c <= 9'b100101110;
				8'b110010: c <= 9'b1011000;
				8'b1101101: c <= 9'b10010000;
				8'b100011: c <= 9'b11011100;
				8'b1110101: c <= 9'b110100001;
				8'b1111101: c <= 9'b11011100;
				8'b101001: c <= 9'b110000011;
				8'b1010010: c <= 9'b110001100;
				8'b1011000: c <= 9'b11101111;
				8'b101110: c <= 9'b110001110;
				8'b1000001: c <= 9'b111111111;
				default: c <= 9'b0;
			endcase
			9'b110111 : case(di)
				8'b1000011: c <= 9'b110001001;
				8'b101000: c <= 9'b10011111;
				8'b111010: c <= 9'b110000101;
				8'b110110: c <= 9'b101110010;
				8'b1100100: c <= 9'b101000101;
				8'b1000000: c <= 9'b110011;
				8'b1110110: c <= 9'b100010111;
				8'b100101: c <= 9'b101101101;
				8'b101111: c <= 9'b101010001;
				8'b100110: c <= 9'b10111000;
				8'b1100011: c <= 9'b10001101;
				8'b1001000: c <= 9'b111110011;
				8'b111000: c <= 9'b11110100;
				8'b110001: c <= 9'b110100010;
				8'b1010111: c <= 9'b101011110;
				8'b1001110: c <= 9'b11110111;
				8'b1101010: c <= 9'b10011011;
				8'b1001001: c <= 9'b11101101;
				8'b1100000: c <= 9'b10000110;
				8'b110111: c <= 9'b1;
				8'b1011101: c <= 9'b11011011;
				8'b1011011: c <= 9'b110101;
				8'b111001: c <= 9'b100101;
				8'b1001010: c <= 9'b101100000;
				8'b110011: c <= 9'b110110000;
				8'b1101100: c <= 9'b111010001;
				8'b1110111: c <= 9'b111001011;
				8'b101011: c <= 9'b1001;
				8'b1101011: c <= 9'b101011110;
				8'b111100: c <= 9'b1101000;
				8'b1000111: c <= 9'b111111101;
				8'b1011111: c <= 9'b1101100;
				8'b1110100: c <= 9'b1011100;
				8'b101101: c <= 9'b11000000;
				8'b1010011: c <= 9'b100001101;
				8'b1100001: c <= 9'b100001110;
				8'b110101: c <= 9'b101101100;
				8'b1000100: c <= 9'b11010001;
				8'b1010001: c <= 9'b100100111;
				8'b1010100: c <= 9'b100000011;
				8'b1100110: c <= 9'b110011110;
				8'b101010: c <= 9'b1011110;
				8'b1011110: c <= 9'b1000100;
				8'b1100111: c <= 9'b111100000;
				8'b1011010: c <= 9'b110011101;
				8'b1000010: c <= 9'b110110010;
				8'b111101: c <= 9'b11101100;
				8'b110000: c <= 9'b100100111;
				8'b111110: c <= 9'b111100111;
				8'b1100010: c <= 9'b1101101;
				8'b1110000: c <= 9'b11011110;
				8'b1101001: c <= 9'b1111000;
				8'b1110011: c <= 9'b110111110;
				8'b1001100: c <= 9'b10110001;
				8'b100001: c <= 9'b101010110;
				8'b1000110: c <= 9'b100111011;
				8'b1110010: c <= 9'b110101101;
				8'b1010000: c <= 9'b110111010;
				8'b1111010: c <= 9'b111000010;
				8'b1010101: c <= 9'b100011111;
				8'b111011: c <= 9'b111000;
				8'b1001101: c <= 9'b11100001;
				8'b111111: c <= 9'b111001011;
				8'b1101110: c <= 9'b111100000;
				8'b1111011: c <= 9'b101001001;
				8'b1001011: c <= 9'b100000110;
				8'b1101111: c <= 9'b10101;
				8'b1101000: c <= 9'b100000111;
				8'b101100: c <= 9'b10100011;
				8'b100100: c <= 9'b101111111;
				8'b1111000: c <= 9'b110101001;
				8'b1000101: c <= 9'b111111111;
				8'b1011001: c <= 9'b110100110;
				8'b110100: c <= 9'b111111101;
				8'b1111001: c <= 9'b111111000;
				8'b1110001: c <= 9'b1001;
				8'b1001111: c <= 9'b100101011;
				8'b1100101: c <= 9'b100;
				8'b1111110: c <= 9'b11111101;
				8'b1111100: c <= 9'b101101110;
				8'b1010110: c <= 9'b11010011;
				8'b110010: c <= 9'b110001111;
				8'b1101101: c <= 9'b1110000;
				8'b100011: c <= 9'b10011111;
				8'b1110101: c <= 9'b101100000;
				8'b1111101: c <= 9'b101010111;
				8'b101001: c <= 9'b11010000;
				8'b1010010: c <= 9'b10001001;
				8'b1011000: c <= 9'b110101101;
				8'b101110: c <= 9'b10000111;
				8'b1000001: c <= 9'b110001;
				default: c <= 9'b0;
			endcase
			9'b101100000 : case(di)
				8'b1000011: c <= 9'b10110001;
				8'b101000: c <= 9'b1011100;
				8'b111010: c <= 9'b11110000;
				8'b110110: c <= 9'b101;
				8'b1100100: c <= 9'b110000;
				8'b1000000: c <= 9'b101110010;
				8'b1110110: c <= 9'b101001011;
				8'b100101: c <= 9'b1000101;
				8'b101111: c <= 9'b110101011;
				8'b100110: c <= 9'b111000101;
				8'b1100011: c <= 9'b10111000;
				8'b1001000: c <= 9'b1011001;
				8'b111000: c <= 9'b100100110;
				8'b110001: c <= 9'b10101010;
				8'b1010111: c <= 9'b111010110;
				8'b1001110: c <= 9'b110100101;
				8'b1101010: c <= 9'b101001111;
				8'b1001001: c <= 9'b100101100;
				8'b1100000: c <= 9'b11011001;
				8'b110111: c <= 9'b101110001;
				8'b1011101: c <= 9'b11111101;
				8'b1011011: c <= 9'b1000010;
				8'b111001: c <= 9'b100011000;
				8'b1001010: c <= 9'b11100111;
				8'b110011: c <= 9'b1111111;
				8'b1101100: c <= 9'b11010001;
				8'b1110111: c <= 9'b111100000;
				8'b101011: c <= 9'b110101110;
				8'b1101011: c <= 9'b11011101;
				8'b111100: c <= 9'b10100110;
				8'b1000111: c <= 9'b100101010;
				8'b1011111: c <= 9'b11000010;
				8'b1110100: c <= 9'b100011011;
				8'b101101: c <= 9'b110110111;
				8'b1010011: c <= 9'b10111110;
				8'b1100001: c <= 9'b1100100;
				8'b110101: c <= 9'b100110100;
				8'b1000100: c <= 9'b100001010;
				8'b1010001: c <= 9'b101001001;
				8'b1010100: c <= 9'b101111001;
				8'b1100110: c <= 9'b111001001;
				8'b101010: c <= 9'b101100010;
				8'b1011110: c <= 9'b11001010;
				8'b1100111: c <= 9'b11000000;
				8'b1011010: c <= 9'b101000101;
				8'b1000010: c <= 9'b100001001;
				8'b111101: c <= 9'b10001011;
				8'b110000: c <= 9'b1110010;
				8'b111110: c <= 9'b1101101;
				8'b1100010: c <= 9'b111100100;
				8'b1110000: c <= 9'b111110011;
				8'b1101001: c <= 9'b111010000;
				8'b1110011: c <= 9'b1101000;
				8'b1001100: c <= 9'b111001001;
				8'b100001: c <= 9'b100001111;
				8'b1000110: c <= 9'b10101101;
				8'b1110010: c <= 9'b11110010;
				8'b1010000: c <= 9'b101111000;
				8'b1111010: c <= 9'b11001110;
				8'b1010101: c <= 9'b1010010;
				8'b111011: c <= 9'b101011110;
				8'b1001101: c <= 9'b110111000;
				8'b111111: c <= 9'b101010011;
				8'b1101110: c <= 9'b10111111;
				8'b1111011: c <= 9'b1100;
				8'b1001011: c <= 9'b11011;
				8'b1101111: c <= 9'b100010011;
				8'b1101000: c <= 9'b111001110;
				8'b101100: c <= 9'b101101001;
				8'b100100: c <= 9'b101001011;
				8'b1111000: c <= 9'b111100;
				8'b1000101: c <= 9'b10100011;
				8'b1011001: c <= 9'b111110001;
				8'b110100: c <= 9'b111000110;
				8'b1111001: c <= 9'b11111110;
				8'b1110001: c <= 9'b110100001;
				8'b1001111: c <= 9'b110001111;
				8'b1100101: c <= 9'b110101010;
				8'b1111110: c <= 9'b10000111;
				8'b1111100: c <= 9'b100000010;
				8'b1010110: c <= 9'b110110011;
				8'b110010: c <= 9'b11001010;
				8'b1101101: c <= 9'b110100100;
				8'b100011: c <= 9'b110011010;
				8'b1110101: c <= 9'b10000;
				8'b1111101: c <= 9'b101000111;
				8'b101001: c <= 9'b10100111;
				8'b1010010: c <= 9'b11100010;
				8'b1011000: c <= 9'b110100100;
				8'b101110: c <= 9'b101100111;
				8'b1000001: c <= 9'b110100110;
				default: c <= 9'b0;
			endcase
			9'b110 : case(di)
				8'b1000011: c <= 9'b111110110;
				8'b101000: c <= 9'b101110101;
				8'b111010: c <= 9'b1001111;
				8'b110110: c <= 9'b10011;
				8'b1100100: c <= 9'b10111;
				8'b1000000: c <= 9'b1011111;
				8'b1110110: c <= 9'b110101110;
				8'b100101: c <= 9'b101101000;
				8'b101111: c <= 9'b11000000;
				8'b100110: c <= 9'b111101000;
				8'b1100011: c <= 9'b10010;
				8'b1001000: c <= 9'b100010111;
				8'b111000: c <= 9'b101110;
				8'b110001: c <= 9'b110100010;
				8'b1010111: c <= 9'b101001011;
				8'b1001110: c <= 9'b110;
				8'b1101010: c <= 9'b101110101;
				8'b1001001: c <= 9'b110001100;
				8'b1100000: c <= 9'b100100110;
				8'b110111: c <= 9'b100011111;
				8'b1011101: c <= 9'b111111101;
				8'b1011011: c <= 9'b110111;
				8'b111001: c <= 9'b101100000;
				8'b1001010: c <= 9'b101100010;
				8'b110011: c <= 9'b100101110;
				8'b1101100: c <= 9'b101010;
				8'b1110111: c <= 9'b101011011;
				8'b101011: c <= 9'b101101000;
				8'b1101011: c <= 9'b100101100;
				8'b111100: c <= 9'b101110100;
				8'b1000111: c <= 9'b100001001;
				8'b1011111: c <= 9'b101010;
				8'b1110100: c <= 9'b1101000;
				8'b101101: c <= 9'b11110110;
				8'b1010011: c <= 9'b110111010;
				8'b1100001: c <= 9'b1101000;
				8'b110101: c <= 9'b101000101;
				8'b1000100: c <= 9'b101000011;
				8'b1010001: c <= 9'b100001100;
				8'b1010100: c <= 9'b10110111;
				8'b1100110: c <= 9'b101110000;
				8'b101010: c <= 9'b10110010;
				8'b1011110: c <= 9'b11110000;
				8'b1100111: c <= 9'b100001100;
				8'b1011010: c <= 9'b100011101;
				8'b1000010: c <= 9'b10111000;
				8'b111101: c <= 9'b10111101;
				8'b110000: c <= 9'b11011100;
				8'b111110: c <= 9'b10000000;
				8'b1100010: c <= 9'b100111110;
				8'b1110000: c <= 9'b10011101;
				8'b1101001: c <= 9'b110110000;
				8'b1110011: c <= 9'b100000111;
				8'b1001100: c <= 9'b110001010;
				8'b100001: c <= 9'b110111111;
				8'b1000110: c <= 9'b111111010;
				8'b1110010: c <= 9'b11111101;
				8'b1010000: c <= 9'b100111111;
				8'b1111010: c <= 9'b10000001;
				8'b1010101: c <= 9'b100010000;
				8'b111011: c <= 9'b111000101;
				8'b1001101: c <= 9'b111111001;
				8'b111111: c <= 9'b111000010;
				8'b1101110: c <= 9'b100110;
				8'b1111011: c <= 9'b101111010;
				8'b1001011: c <= 9'b100000101;
				8'b1101111: c <= 9'b101101011;
				8'b1101000: c <= 9'b100000100;
				8'b101100: c <= 9'b101101010;
				8'b100100: c <= 9'b10001000;
				8'b1111000: c <= 9'b111101;
				8'b1000101: c <= 9'b10110;
				8'b1011001: c <= 9'b111110011;
				8'b110100: c <= 9'b10001110;
				8'b1111001: c <= 9'b111011110;
				8'b1110001: c <= 9'b11001110;
				8'b1001111: c <= 9'b111001111;
				8'b1100101: c <= 9'b100001111;
				8'b1111110: c <= 9'b11001000;
				8'b1111100: c <= 9'b111000011;
				8'b1010110: c <= 9'b10111000;
				8'b110010: c <= 9'b111000101;
				8'b1101101: c <= 9'b11111101;
				8'b100011: c <= 9'b101000111;
				8'b1110101: c <= 9'b11101011;
				8'b1111101: c <= 9'b1110100;
				8'b101001: c <= 9'b10000111;
				8'b1010010: c <= 9'b100111000;
				8'b1011000: c <= 9'b111010110;
				8'b101110: c <= 9'b10010100;
				8'b1000001: c <= 9'b1110111;
				default: c <= 9'b0;
			endcase
			9'b1001011 : case(di)
				8'b1000011: c <= 9'b10110;
				8'b101000: c <= 9'b101010101;
				8'b111010: c <= 9'b10011001;
				8'b110110: c <= 9'b111101010;
				8'b1100100: c <= 9'b10100000;
				8'b1000000: c <= 9'b1101101;
				8'b1110110: c <= 9'b10010110;
				8'b100101: c <= 9'b10101000;
				8'b101111: c <= 9'b1111;
				8'b100110: c <= 9'b10111011;
				8'b1100011: c <= 9'b11001110;
				8'b1001000: c <= 9'b11111110;
				8'b111000: c <= 9'b1110111;
				8'b110001: c <= 9'b1000011;
				8'b1010111: c <= 9'b1001100;
				8'b1001110: c <= 9'b100000011;
				8'b1101010: c <= 9'b101001110;
				8'b1001001: c <= 9'b11011001;
				8'b1100000: c <= 9'b1001010;
				8'b110111: c <= 9'b101110100;
				8'b1011101: c <= 9'b110111000;
				8'b1011011: c <= 9'b101101010;
				8'b111001: c <= 9'b101011;
				8'b1001010: c <= 9'b110111;
				8'b110011: c <= 9'b110100110;
				8'b1101100: c <= 9'b10001111;
				8'b1110111: c <= 9'b110100101;
				8'b101011: c <= 9'b10111110;
				8'b1101011: c <= 9'b10100110;
				8'b111100: c <= 9'b111011011;
				8'b1000111: c <= 9'b11001001;
				8'b1011111: c <= 9'b11100111;
				8'b1110100: c <= 9'b100100000;
				8'b101101: c <= 9'b11010000;
				8'b1010011: c <= 9'b101010;
				8'b1100001: c <= 9'b100100010;
				8'b110101: c <= 9'b11111101;
				8'b1000100: c <= 9'b1111010;
				8'b1010001: c <= 9'b110011101;
				8'b1010100: c <= 9'b1110111;
				8'b1100110: c <= 9'b11101011;
				8'b101010: c <= 9'b101001011;
				8'b1011110: c <= 9'b101011010;
				8'b1100111: c <= 9'b1001001;
				8'b1011010: c <= 9'b101101000;
				8'b1000010: c <= 9'b110100101;
				8'b111101: c <= 9'b11111100;
				8'b110000: c <= 9'b10001011;
				8'b111110: c <= 9'b111110101;
				8'b1100010: c <= 9'b11001000;
				8'b1110000: c <= 9'b1101110;
				8'b1101001: c <= 9'b111000011;
				8'b1110011: c <= 9'b10111000;
				8'b1001100: c <= 9'b1110111;
				8'b100001: c <= 9'b111111011;
				8'b1000110: c <= 9'b11111101;
				8'b1110010: c <= 9'b111010100;
				8'b1010000: c <= 9'b1001001;
				8'b1111010: c <= 9'b100001111;
				8'b1010101: c <= 9'b10001011;
				8'b111011: c <= 9'b100001;
				8'b1001101: c <= 9'b10010100;
				8'b111111: c <= 9'b111010111;
				8'b1101110: c <= 9'b111010111;
				8'b1111011: c <= 9'b111110000;
				8'b1001011: c <= 9'b1100110;
				8'b1101111: c <= 9'b1101110;
				8'b1101000: c <= 9'b110011;
				8'b101100: c <= 9'b111110101;
				8'b100100: c <= 9'b110111001;
				8'b1111000: c <= 9'b11110110;
				8'b1000101: c <= 9'b100011;
				8'b1011001: c <= 9'b101111010;
				8'b110100: c <= 9'b100100110;
				8'b1111001: c <= 9'b10000111;
				8'b1110001: c <= 9'b11011101;
				8'b1001111: c <= 9'b10001010;
				8'b1100101: c <= 9'b100110111;
				8'b1111110: c <= 9'b111011011;
				8'b1111100: c <= 9'b1110100;
				8'b1010110: c <= 9'b1111001;
				8'b110010: c <= 9'b100100110;
				8'b1101101: c <= 9'b10100000;
				8'b100011: c <= 9'b10011100;
				8'b1110101: c <= 9'b101000010;
				8'b1111101: c <= 9'b10000001;
				8'b101001: c <= 9'b110011000;
				8'b1010010: c <= 9'b1101000;
				8'b1011000: c <= 9'b101100000;
				8'b101110: c <= 9'b10000110;
				8'b1000001: c <= 9'b101001111;
				default: c <= 9'b0;
			endcase
			9'b1000101 : case(di)
				8'b1000011: c <= 9'b101110100;
				8'b101000: c <= 9'b101010;
				8'b111010: c <= 9'b100011100;
				8'b110110: c <= 9'b110010111;
				8'b1100100: c <= 9'b1000011;
				8'b1000000: c <= 9'b100000001;
				8'b1110110: c <= 9'b10000;
				8'b100101: c <= 9'b1100001;
				8'b101111: c <= 9'b111010;
				8'b100110: c <= 9'b110100;
				8'b1100011: c <= 9'b100010011;
				8'b1001000: c <= 9'b10001110;
				8'b111000: c <= 9'b110111111;
				8'b110001: c <= 9'b110100011;
				8'b1010111: c <= 9'b110111;
				8'b1001110: c <= 9'b111100011;
				8'b1101010: c <= 9'b100100101;
				8'b1001001: c <= 9'b111100100;
				8'b1100000: c <= 9'b101101111;
				8'b110111: c <= 9'b10100;
				8'b1011101: c <= 9'b100110010;
				8'b1011011: c <= 9'b111;
				8'b111001: c <= 9'b101110001;
				8'b1001010: c <= 9'b110111010;
				8'b110011: c <= 9'b110100111;
				8'b1101100: c <= 9'b11000001;
				8'b1110111: c <= 9'b111001011;
				8'b101011: c <= 9'b1101111;
				8'b1101011: c <= 9'b11010101;
				8'b111100: c <= 9'b111001100;
				8'b1000111: c <= 9'b111001;
				8'b1011111: c <= 9'b10011010;
				8'b1110100: c <= 9'b100011001;
				8'b101101: c <= 9'b111101111;
				8'b1010011: c <= 9'b10001110;
				8'b1100001: c <= 9'b1111110;
				8'b110101: c <= 9'b1010010;
				8'b1000100: c <= 9'b1000110;
				8'b1010001: c <= 9'b100100111;
				8'b1010100: c <= 9'b11111010;
				8'b1100110: c <= 9'b10000010;
				8'b101010: c <= 9'b100111110;
				8'b1011110: c <= 9'b11011101;
				8'b1100111: c <= 9'b111001110;
				8'b1011010: c <= 9'b101010110;
				8'b1000010: c <= 9'b11101011;
				8'b111101: c <= 9'b1001100;
				8'b110000: c <= 9'b111101010;
				8'b111110: c <= 9'b111111101;
				8'b1100010: c <= 9'b10110110;
				8'b1110000: c <= 9'b110101110;
				8'b1101001: c <= 9'b100111;
				8'b1110011: c <= 9'b100000000;
				8'b1001100: c <= 9'b101110010;
				8'b100001: c <= 9'b100010100;
				8'b1000110: c <= 9'b101000011;
				8'b1110010: c <= 9'b11001111;
				8'b1010000: c <= 9'b11010100;
				8'b1111010: c <= 9'b111101110;
				8'b1010101: c <= 9'b111001110;
				8'b111011: c <= 9'b111000100;
				8'b1001101: c <= 9'b110100000;
				8'b111111: c <= 9'b100100000;
				8'b1101110: c <= 9'b101000001;
				8'b1111011: c <= 9'b110011111;
				8'b1001011: c <= 9'b101011;
				8'b1101111: c <= 9'b1010010;
				8'b1101000: c <= 9'b101100101;
				8'b101100: c <= 9'b111000100;
				8'b100100: c <= 9'b111010100;
				8'b1111000: c <= 9'b10010111;
				8'b1000101: c <= 9'b101000100;
				8'b1011001: c <= 9'b11111;
				8'b110100: c <= 9'b101110100;
				8'b1111001: c <= 9'b11011010;
				8'b1110001: c <= 9'b11100000;
				8'b1001111: c <= 9'b100110110;
				8'b1100101: c <= 9'b101110101;
				8'b1111110: c <= 9'b10000000;
				8'b1111100: c <= 9'b111111011;
				8'b1010110: c <= 9'b100111;
				8'b110010: c <= 9'b110001;
				8'b1101101: c <= 9'b111101;
				8'b100011: c <= 9'b11111;
				8'b1110101: c <= 9'b10100100;
				8'b1111101: c <= 9'b10100010;
				8'b101001: c <= 9'b1001;
				8'b1010010: c <= 9'b111011001;
				8'b1011000: c <= 9'b111000011;
				8'b101110: c <= 9'b101011101;
				8'b1000001: c <= 9'b111001011;
				default: c <= 9'b0;
			endcase
			9'b1001 : case(di)
				8'b1000011: c <= 9'b11101100;
				8'b101000: c <= 9'b100111101;
				8'b111010: c <= 9'b101101000;
				8'b110110: c <= 9'b11100010;
				8'b1100100: c <= 9'b110110111;
				8'b1000000: c <= 9'b110110011;
				8'b1110110: c <= 9'b1000010;
				8'b100101: c <= 9'b100000000;
				8'b101111: c <= 9'b110011;
				8'b100110: c <= 9'b10111001;
				8'b1100011: c <= 9'b101010111;
				8'b1001000: c <= 9'b10000101;
				8'b111000: c <= 9'b110011111;
				8'b110001: c <= 9'b1101111;
				8'b1010111: c <= 9'b111111011;
				8'b1001110: c <= 9'b101000011;
				8'b1101010: c <= 9'b11010101;
				8'b1001001: c <= 9'b11111101;
				8'b1100000: c <= 9'b111000000;
				8'b110111: c <= 9'b110010011;
				8'b1011101: c <= 9'b100111100;
				8'b1011011: c <= 9'b111001111;
				8'b111001: c <= 9'b111011001;
				8'b1001010: c <= 9'b101000011;
				8'b110011: c <= 9'b11001;
				8'b1101100: c <= 9'b110100;
				8'b1110111: c <= 9'b110101101;
				8'b101011: c <= 9'b11110101;
				8'b1101011: c <= 9'b1011100;
				8'b111100: c <= 9'b1100011;
				8'b1000111: c <= 9'b111110000;
				8'b1011111: c <= 9'b1001101;
				8'b1110100: c <= 9'b100001;
				8'b101101: c <= 9'b101000101;
				8'b1010011: c <= 9'b101101111;
				8'b1100001: c <= 9'b101000;
				8'b110101: c <= 9'b1011010;
				8'b1000100: c <= 9'b111111110;
				8'b1010001: c <= 9'b100011101;
				8'b1010100: c <= 9'b110100000;
				8'b1100110: c <= 9'b110100110;
				8'b101010: c <= 9'b11000110;
				8'b1011110: c <= 9'b10101010;
				8'b1100111: c <= 9'b111111001;
				8'b1011010: c <= 9'b110111011;
				8'b1000010: c <= 9'b101100111;
				8'b111101: c <= 9'b110001010;
				8'b110000: c <= 9'b110101101;
				8'b111110: c <= 9'b1001000;
				8'b1100010: c <= 9'b111001101;
				8'b1110000: c <= 9'b111001111;
				8'b1101001: c <= 9'b10111000;
				8'b1110011: c <= 9'b111010010;
				8'b1001100: c <= 9'b111000111;
				8'b100001: c <= 9'b110000010;
				8'b1000110: c <= 9'b111101000;
				8'b1110010: c <= 9'b111111101;
				8'b1010000: c <= 9'b100011011;
				8'b1111010: c <= 9'b101100100;
				8'b1010101: c <= 9'b101010101;
				8'b111011: c <= 9'b1100011;
				8'b1001101: c <= 9'b111100100;
				8'b111111: c <= 9'b101110100;
				8'b1101110: c <= 9'b11001;
				8'b1111011: c <= 9'b10010101;
				8'b1001011: c <= 9'b11100110;
				8'b1101111: c <= 9'b11100;
				8'b1101000: c <= 9'b101101001;
				8'b101100: c <= 9'b1001110;
				8'b100100: c <= 9'b10110101;
				8'b1111000: c <= 9'b10000;
				8'b1000101: c <= 9'b101;
				8'b1011001: c <= 9'b10100101;
				8'b110100: c <= 9'b10101001;
				8'b1111001: c <= 9'b100111111;
				8'b1110001: c <= 9'b101001001;
				8'b1001111: c <= 9'b11010;
				8'b1100101: c <= 9'b111010100;
				8'b1111110: c <= 9'b1001011;
				8'b1111100: c <= 9'b101100000;
				8'b1010110: c <= 9'b11110110;
				8'b110010: c <= 9'b101100101;
				8'b1101101: c <= 9'b100011001;
				8'b100011: c <= 9'b100100011;
				8'b1110101: c <= 9'b101110101;
				8'b1111101: c <= 9'b101110100;
				8'b101001: c <= 9'b111100010;
				8'b1010010: c <= 9'b100110100;
				8'b1011000: c <= 9'b111101101;
				8'b101110: c <= 9'b10000001;
				8'b1000001: c <= 9'b10101010;
				default: c <= 9'b0;
			endcase
			9'b10110011 : case(di)
				8'b1000011: c <= 9'b10001110;
				8'b101000: c <= 9'b100100110;
				8'b111010: c <= 9'b11010001;
				8'b110110: c <= 9'b111001011;
				8'b1100100: c <= 9'b101100100;
				8'b1000000: c <= 9'b111010000;
				8'b1110110: c <= 9'b11001001;
				8'b100101: c <= 9'b101111000;
				8'b101111: c <= 9'b11100000;
				8'b100110: c <= 9'b111000100;
				8'b1100011: c <= 9'b1001011;
				8'b1001000: c <= 9'b101100000;
				8'b111000: c <= 9'b10110;
				8'b110001: c <= 9'b110000010;
				8'b1010111: c <= 9'b1010010;
				8'b1001110: c <= 9'b1101000;
				8'b1101010: c <= 9'b11100010;
				8'b1001001: c <= 9'b100000101;
				8'b1100000: c <= 9'b1001;
				8'b110111: c <= 9'b1101100;
				8'b1011101: c <= 9'b11100011;
				8'b1011011: c <= 9'b111000011;
				8'b111001: c <= 9'b100;
				8'b1001010: c <= 9'b1000000;
				8'b110011: c <= 9'b10010101;
				8'b1101100: c <= 9'b1100110;
				8'b1110111: c <= 9'b101101000;
				8'b101011: c <= 9'b110011110;
				8'b1101011: c <= 9'b100111010;
				8'b111100: c <= 9'b100110111;
				8'b1000111: c <= 9'b1111011;
				8'b1011111: c <= 9'b10000110;
				8'b1110100: c <= 9'b111110101;
				8'b101101: c <= 9'b101110101;
				8'b1010011: c <= 9'b101011101;
				8'b1100001: c <= 9'b111101;
				8'b110101: c <= 9'b110110000;
				8'b1000100: c <= 9'b1111000;
				8'b1010001: c <= 9'b100110011;
				8'b1010100: c <= 9'b1111100;
				8'b1100110: c <= 9'b100101111;
				8'b101010: c <= 9'b101100100;
				8'b1011110: c <= 9'b10010011;
				8'b1100111: c <= 9'b101101011;
				8'b1011010: c <= 9'b101110010;
				8'b1000010: c <= 9'b101011111;
				8'b111101: c <= 9'b101010;
				8'b110000: c <= 9'b10000010;
				8'b111110: c <= 9'b100101101;
				8'b1100010: c <= 9'b100101;
				8'b1110000: c <= 9'b1110111;
				8'b1101001: c <= 9'b110000001;
				8'b1110011: c <= 9'b110110000;
				8'b1001100: c <= 9'b100110111;
				8'b100001: c <= 9'b100111001;
				8'b1000110: c <= 9'b111;
				8'b1110010: c <= 9'b11111010;
				8'b1010000: c <= 9'b101100000;
				8'b1111010: c <= 9'b10000011;
				8'b1010101: c <= 9'b11100101;
				8'b111011: c <= 9'b111100001;
				8'b1001101: c <= 9'b1101000;
				8'b111111: c <= 9'b10111011;
				8'b1101110: c <= 9'b110101110;
				8'b1111011: c <= 9'b11011101;
				8'b1001011: c <= 9'b101101010;
				8'b1101111: c <= 9'b110010001;
				8'b1101000: c <= 9'b101000;
				8'b101100: c <= 9'b10101110;
				8'b100100: c <= 9'b110101001;
				8'b1111000: c <= 9'b100101001;
				8'b1000101: c <= 9'b111001100;
				8'b1011001: c <= 9'b110011100;
				8'b110100: c <= 9'b1110011;
				8'b1111001: c <= 9'b111001;
				8'b1110001: c <= 9'b100000100;
				8'b1001111: c <= 9'b11100111;
				8'b1100101: c <= 9'b111010;
				8'b1111110: c <= 9'b10101000;
				8'b1111100: c <= 9'b10;
				8'b1010110: c <= 9'b100001111;
				8'b110010: c <= 9'b101110111;
				8'b1101101: c <= 9'b1101111;
				8'b100011: c <= 9'b10000011;
				8'b1110101: c <= 9'b110110101;
				8'b1111101: c <= 9'b110110100;
				8'b101001: c <= 9'b101111010;
				8'b1010010: c <= 9'b11000110;
				8'b1011000: c <= 9'b110000111;
				8'b101110: c <= 9'b110000001;
				8'b1000001: c <= 9'b111010110;
				default: c <= 9'b0;
			endcase
			9'b110100011 : case(di)
				8'b1000011: c <= 9'b111001111;
				8'b101000: c <= 9'b10101001;
				8'b111010: c <= 9'b111101100;
				8'b110110: c <= 9'b1100111;
				8'b1100100: c <= 9'b11100010;
				8'b1000000: c <= 9'b1111101;
				8'b1110110: c <= 9'b100011101;
				8'b100101: c <= 9'b1100000;
				8'b101111: c <= 9'b101110101;
				8'b100110: c <= 9'b100111010;
				8'b1100011: c <= 9'b1100110;
				8'b1001000: c <= 9'b111011;
				8'b111000: c <= 9'b101000011;
				8'b110001: c <= 9'b10011001;
				8'b1010111: c <= 9'b10111000;
				8'b1001110: c <= 9'b110101011;
				8'b1101010: c <= 9'b110101;
				8'b1001001: c <= 9'b110101010;
				8'b1100000: c <= 9'b10010011;
				8'b110111: c <= 9'b110101101;
				8'b1011101: c <= 9'b10100;
				8'b1011011: c <= 9'b1101001;
				8'b111001: c <= 9'b1100101;
				8'b1001010: c <= 9'b1010111;
				8'b110011: c <= 9'b101110101;
				8'b1101100: c <= 9'b100010110;
				8'b1110111: c <= 9'b111101;
				8'b101011: c <= 9'b111011111;
				8'b1101011: c <= 9'b111000111;
				8'b111100: c <= 9'b100101001;
				8'b1000111: c <= 9'b110011101;
				8'b1011111: c <= 9'b110011001;
				8'b1110100: c <= 9'b110010110;
				8'b101101: c <= 9'b101100010;
				8'b1010011: c <= 9'b100000110;
				8'b1100001: c <= 9'b101001011;
				8'b110101: c <= 9'b1111000;
				8'b1000100: c <= 9'b100001010;
				8'b1010001: c <= 9'b1100010;
				8'b1010100: c <= 9'b10100110;
				8'b1100110: c <= 9'b11111010;
				8'b101010: c <= 9'b100001001;
				8'b1011110: c <= 9'b110001101;
				8'b1100111: c <= 9'b10101;
				8'b1011010: c <= 9'b110000011;
				8'b1000010: c <= 9'b111101010;
				8'b111101: c <= 9'b1010001;
				8'b110000: c <= 9'b1110010;
				8'b111110: c <= 9'b10111010;
				8'b1100010: c <= 9'b101101010;
				8'b1110000: c <= 9'b11001;
				8'b1101001: c <= 9'b1011010;
				8'b1110011: c <= 9'b11000111;
				8'b1001100: c <= 9'b1001;
				8'b100001: c <= 9'b1111100;
				8'b1000110: c <= 9'b11010101;
				8'b1110010: c <= 9'b101010101;
				8'b1010000: c <= 9'b111000010;
				8'b1111010: c <= 9'b11001010;
				8'b1010101: c <= 9'b10101110;
				8'b111011: c <= 9'b110100010;
				8'b1001101: c <= 9'b10111110;
				8'b111111: c <= 9'b110001011;
				8'b1101110: c <= 9'b1110111;
				8'b1111011: c <= 9'b1011010;
				8'b1001011: c <= 9'b111001100;
				8'b1101111: c <= 9'b1111100;
				8'b1101000: c <= 9'b1001000;
				8'b101100: c <= 9'b111;
				8'b100100: c <= 9'b110111100;
				8'b1111000: c <= 9'b101101101;
				8'b1000101: c <= 9'b111000010;
				8'b1011001: c <= 9'b11101001;
				8'b110100: c <= 9'b101101101;
				8'b1111001: c <= 9'b100000110;
				8'b1110001: c <= 9'b111011110;
				8'b1001111: c <= 9'b111011010;
				8'b1100101: c <= 9'b1001010;
				8'b1111110: c <= 9'b110001000;
				8'b1111100: c <= 9'b101001001;
				8'b1010110: c <= 9'b110101011;
				8'b110010: c <= 9'b100010001;
				8'b1101101: c <= 9'b111000010;
				8'b100011: c <= 9'b111;
				8'b1110101: c <= 9'b11001;
				8'b1111101: c <= 9'b1001100;
				8'b101001: c <= 9'b10101011;
				8'b1010010: c <= 9'b10101010;
				8'b1011000: c <= 9'b100111101;
				8'b101110: c <= 9'b111111010;
				8'b1000001: c <= 9'b111111000;
				default: c <= 9'b0;
			endcase
			9'b10111 : case(di)
				8'b1000011: c <= 9'b10011111;
				8'b101000: c <= 9'b110011;
				8'b111010: c <= 9'b10001000;
				8'b110110: c <= 9'b100100001;
				8'b1100100: c <= 9'b100001100;
				8'b1000000: c <= 9'b10110101;
				8'b1110110: c <= 9'b110100;
				8'b100101: c <= 9'b111001000;
				8'b101111: c <= 9'b1100111;
				8'b100110: c <= 9'b101101111;
				8'b1100011: c <= 9'b100100111;
				8'b1001000: c <= 9'b1111011;
				8'b111000: c <= 9'b100011011;
				8'b110001: c <= 9'b111101110;
				8'b1010111: c <= 9'b111011111;
				8'b1001110: c <= 9'b100010101;
				8'b1101010: c <= 9'b111101100;
				8'b1001001: c <= 9'b10100011;
				8'b1100000: c <= 9'b11001111;
				8'b110111: c <= 9'b1011110;
				8'b1011101: c <= 9'b100;
				8'b1011011: c <= 9'b10100100;
				8'b111001: c <= 9'b1100011;
				8'b1001010: c <= 9'b11110000;
				8'b110011: c <= 9'b111001111;
				8'b1101100: c <= 9'b10101011;
				8'b1110111: c <= 9'b11000000;
				8'b101011: c <= 9'b1100100;
				8'b1101011: c <= 9'b10000;
				8'b111100: c <= 9'b101;
				8'b1000111: c <= 9'b1000011;
				8'b1011111: c <= 9'b110010;
				8'b1110100: c <= 9'b101011111;
				8'b101101: c <= 9'b110101001;
				8'b1010011: c <= 9'b101001011;
				8'b1100001: c <= 9'b101101001;
				8'b110101: c <= 9'b1001;
				8'b1000100: c <= 9'b110111001;
				8'b1010001: c <= 9'b1000;
				8'b1010100: c <= 9'b11110000;
				8'b1100110: c <= 9'b111111011;
				8'b101010: c <= 9'b11100100;
				8'b1011110: c <= 9'b111001010;
				8'b1100111: c <= 9'b10000000;
				8'b1011010: c <= 9'b1010000;
				8'b1000010: c <= 9'b11101101;
				8'b111101: c <= 9'b111111011;
				8'b110000: c <= 9'b1100000;
				8'b111110: c <= 9'b101011111;
				8'b1100010: c <= 9'b110000010;
				8'b1110000: c <= 9'b100100010;
				8'b1101001: c <= 9'b100010000;
				8'b1110011: c <= 9'b10100111;
				8'b1001100: c <= 9'b10100111;
				8'b100001: c <= 9'b11000110;
				8'b1000110: c <= 9'b11010111;
				8'b1110010: c <= 9'b101000111;
				8'b1010000: c <= 9'b10001010;
				8'b1111010: c <= 9'b110001000;
				8'b1010101: c <= 9'b101001100;
				8'b111011: c <= 9'b11110;
				8'b1001101: c <= 9'b101110000;
				8'b111111: c <= 9'b100011000;
				8'b1101110: c <= 9'b111101110;
				8'b1111011: c <= 9'b10111100;
				8'b1001011: c <= 9'b101110111;
				8'b1101111: c <= 9'b1011011;
				8'b1101000: c <= 9'b1001101;
				8'b101100: c <= 9'b10101010;
				8'b100100: c <= 9'b110100010;
				8'b1111000: c <= 9'b111011111;
				8'b1000101: c <= 9'b11110001;
				8'b1011001: c <= 9'b111001101;
				8'b110100: c <= 9'b10001101;
				8'b1111001: c <= 9'b110011010;
				8'b1110001: c <= 9'b10111111;
				8'b1001111: c <= 9'b110110110;
				8'b1100101: c <= 9'b100001110;
				8'b1111110: c <= 9'b101101;
				8'b1111100: c <= 9'b10110111;
				8'b1010110: c <= 9'b110101011;
				8'b110010: c <= 9'b1110010;
				8'b1101101: c <= 9'b1111;
				8'b100011: c <= 9'b11010;
				8'b1110101: c <= 9'b101000110;
				8'b1111101: c <= 9'b10010011;
				8'b101001: c <= 9'b100001110;
				8'b1010010: c <= 9'b1101100;
				8'b1011000: c <= 9'b110010011;
				8'b101110: c <= 9'b11000100;
				8'b1000001: c <= 9'b10100111;
				default: c <= 9'b0;
			endcase
			9'b11000011 : case(di)
				8'b1000011: c <= 9'b110110000;
				8'b101000: c <= 9'b10000110;
				8'b111010: c <= 9'b101100;
				8'b110110: c <= 9'b11011000;
				8'b1100100: c <= 9'b10111000;
				8'b1000000: c <= 9'b11000001;
				8'b1110110: c <= 9'b101000110;
				8'b100101: c <= 9'b111000011;
				8'b101111: c <= 9'b1110;
				8'b100110: c <= 9'b11;
				8'b1100011: c <= 9'b10010110;
				8'b1001000: c <= 9'b1001011;
				8'b111000: c <= 9'b111100111;
				8'b110001: c <= 9'b100001100;
				8'b1010111: c <= 9'b101011011;
				8'b1001110: c <= 9'b110111001;
				8'b1101010: c <= 9'b110001100;
				8'b1001001: c <= 9'b100110010;
				8'b1100000: c <= 9'b111110011;
				8'b110111: c <= 9'b111110001;
				8'b1011101: c <= 9'b111000000;
				8'b1011011: c <= 9'b101100011;
				8'b111001: c <= 9'b110001110;
				8'b1001010: c <= 9'b10011011;
				8'b110011: c <= 9'b1010101;
				8'b1101100: c <= 9'b100010;
				8'b1110111: c <= 9'b110110110;
				8'b101011: c <= 9'b10011;
				8'b1101011: c <= 9'b111011011;
				8'b111100: c <= 9'b111101010;
				8'b1000111: c <= 9'b10010111;
				8'b1011111: c <= 9'b11010011;
				8'b1110100: c <= 9'b101011101;
				8'b101101: c <= 9'b11110;
				8'b1010011: c <= 9'b11111110;
				8'b1100001: c <= 9'b101001;
				8'b110101: c <= 9'b101001011;
				8'b1000100: c <= 9'b11000100;
				8'b1010001: c <= 9'b111011001;
				8'b1010100: c <= 9'b1001000;
				8'b1100110: c <= 9'b11010001;
				8'b101010: c <= 9'b110001100;
				8'b1011110: c <= 9'b1101101;
				8'b1100111: c <= 9'b101011111;
				8'b1011010: c <= 9'b1100011;
				8'b1000010: c <= 9'b11110111;
				8'b111101: c <= 9'b111000011;
				8'b110000: c <= 9'b111101100;
				8'b111110: c <= 9'b10111100;
				8'b1100010: c <= 9'b101101000;
				8'b1110000: c <= 9'b10011100;
				8'b1101001: c <= 9'b100100111;
				8'b1110011: c <= 9'b100010000;
				8'b1001100: c <= 9'b101110101;
				8'b100001: c <= 9'b111111010;
				8'b1000110: c <= 9'b110011101;
				8'b1110010: c <= 9'b11100;
				8'b1010000: c <= 9'b10000101;
				8'b1111010: c <= 9'b1011100;
				8'b1010101: c <= 9'b11110001;
				8'b111011: c <= 9'b101100111;
				8'b1001101: c <= 9'b10101000;
				8'b111111: c <= 9'b100001001;
				8'b1101110: c <= 9'b110011;
				8'b1111011: c <= 9'b110100001;
				8'b1001011: c <= 9'b11000000;
				8'b1101111: c <= 9'b11011100;
				8'b1101000: c <= 9'b1111000;
				8'b101100: c <= 9'b101011;
				8'b100100: c <= 9'b100111010;
				8'b1111000: c <= 9'b110000011;
				8'b1000101: c <= 9'b11001011;
				8'b1011001: c <= 9'b10100100;
				8'b110100: c <= 9'b10010000;
				8'b1111001: c <= 9'b11110000;
				8'b1110001: c <= 9'b110111110;
				8'b1001111: c <= 9'b101100001;
				8'b1100101: c <= 9'b101101101;
				8'b1111110: c <= 9'b110111111;
				8'b1111100: c <= 9'b11111;
				8'b1010110: c <= 9'b11000000;
				8'b110010: c <= 9'b111100001;
				8'b1101101: c <= 9'b11100101;
				8'b100011: c <= 9'b101100010;
				8'b1110101: c <= 9'b1000100;
				8'b1111101: c <= 9'b100100;
				8'b101001: c <= 9'b111111111;
				8'b1010010: c <= 9'b111000111;
				8'b1011000: c <= 9'b10111000;
				8'b101110: c <= 9'b1000111;
				8'b1000001: c <= 9'b11001111;
				default: c <= 9'b0;
			endcase
			9'b100111111 : case(di)
				8'b1000011: c <= 9'b110010;
				8'b101000: c <= 9'b1011;
				8'b111010: c <= 9'b100101;
				8'b110110: c <= 9'b110001110;
				8'b1100100: c <= 9'b100001010;
				8'b1000000: c <= 9'b110011001;
				8'b1110110: c <= 9'b110110000;
				8'b100101: c <= 9'b101001110;
				8'b101111: c <= 9'b1111111;
				8'b100110: c <= 9'b10011101;
				8'b1100011: c <= 9'b101011111;
				8'b1001000: c <= 9'b101011110;
				8'b111000: c <= 9'b100011101;
				8'b110001: c <= 9'b11111101;
				8'b1010111: c <= 9'b11000010;
				8'b1001110: c <= 9'b11110000;
				8'b1101010: c <= 9'b111010110;
				8'b1001001: c <= 9'b101101001;
				8'b1100000: c <= 9'b101110001;
				8'b110111: c <= 9'b110101010;
				8'b1011101: c <= 9'b101000011;
				8'b1011011: c <= 9'b1000111;
				8'b111001: c <= 9'b10100;
				8'b1001010: c <= 9'b100001111;
				8'b110011: c <= 9'b100111111;
				8'b1101100: c <= 9'b110011001;
				8'b1110111: c <= 9'b110111;
				8'b101011: c <= 9'b10001000;
				8'b1101011: c <= 9'b1000000;
				8'b111100: c <= 9'b10001011;
				8'b1000111: c <= 9'b101101010;
				8'b1011111: c <= 9'b11100111;
				8'b1110100: c <= 9'b10010001;
				8'b101101: c <= 9'b101110011;
				8'b1010011: c <= 9'b111011111;
				8'b1100001: c <= 9'b111010001;
				8'b110101: c <= 9'b100100011;
				8'b1000100: c <= 9'b101000001;
				8'b1010001: c <= 9'b111000110;
				8'b1010100: c <= 9'b110000101;
				8'b1100110: c <= 9'b11011000;
				8'b101010: c <= 9'b100010011;
				8'b1011110: c <= 9'b111111;
				8'b1100111: c <= 9'b10000011;
				8'b1011010: c <= 9'b101101010;
				8'b1000010: c <= 9'b10000001;
				8'b111101: c <= 9'b110110100;
				8'b110000: c <= 9'b110000110;
				8'b111110: c <= 9'b111111010;
				8'b1100010: c <= 9'b1111000;
				8'b1110000: c <= 9'b101101011;
				8'b1101001: c <= 9'b10001110;
				8'b1110011: c <= 9'b11000100;
				8'b1001100: c <= 9'b101001100;
				8'b100001: c <= 9'b11111000;
				8'b1000110: c <= 9'b111100000;
				8'b1110010: c <= 9'b110111010;
				8'b1010000: c <= 9'b101010001;
				8'b1111010: c <= 9'b10100100;
				8'b1010101: c <= 9'b100010110;
				8'b111011: c <= 9'b111101111;
				8'b1001101: c <= 9'b11000111;
				8'b111111: c <= 9'b101111110;
				8'b1101110: c <= 9'b101111000;
				8'b1111011: c <= 9'b11010101;
				8'b1001011: c <= 9'b110100011;
				8'b1101111: c <= 9'b110000000;
				8'b1101000: c <= 9'b1000;
				8'b101100: c <= 9'b1111000;
				8'b100100: c <= 9'b11011100;
				8'b1111000: c <= 9'b100110011;
				8'b1000101: c <= 9'b11101000;
				8'b1011001: c <= 9'b111111110;
				8'b110100: c <= 9'b111011111;
				8'b1111001: c <= 9'b111001110;
				8'b1110001: c <= 9'b10;
				8'b1001111: c <= 9'b11101011;
				8'b1100101: c <= 9'b1111101;
				8'b1111110: c <= 9'b101011000;
				8'b1111100: c <= 9'b11010111;
				8'b1010110: c <= 9'b11000;
				8'b110010: c <= 9'b11100101;
				8'b1101101: c <= 9'b1001100;
				8'b100011: c <= 9'b100011100;
				8'b1110101: c <= 9'b100000111;
				8'b1111101: c <= 9'b101100011;
				8'b101001: c <= 9'b10010;
				8'b1010010: c <= 9'b111001001;
				8'b1011000: c <= 9'b111101010;
				8'b101110: c <= 9'b1011011;
				8'b1000001: c <= 9'b100101101;
				default: c <= 9'b0;
			endcase
			9'b10100100 : case(di)
				8'b1000011: c <= 9'b1111101;
				8'b101000: c <= 9'b10000101;
				8'b111010: c <= 9'b1111001;
				8'b110110: c <= 9'b100011011;
				8'b1100100: c <= 9'b100010110;
				8'b1000000: c <= 9'b10011000;
				8'b1110110: c <= 9'b111001111;
				8'b100101: c <= 9'b11000001;
				8'b101111: c <= 9'b101011;
				8'b100110: c <= 9'b11000000;
				8'b1100011: c <= 9'b100110011;
				8'b1001000: c <= 9'b110010010;
				8'b111000: c <= 9'b111101000;
				8'b110001: c <= 9'b11010111;
				8'b1010111: c <= 9'b101110000;
				8'b1001110: c <= 9'b11010001;
				8'b1101010: c <= 9'b11011100;
				8'b1001001: c <= 9'b111101111;
				8'b1100000: c <= 9'b100111101;
				8'b110111: c <= 9'b101011111;
				8'b1011101: c <= 9'b110011;
				8'b1011011: c <= 9'b10011100;
				8'b111001: c <= 9'b101110101;
				8'b1001010: c <= 9'b11010111;
				8'b110011: c <= 9'b10011;
				8'b1101100: c <= 9'b100110101;
				8'b1110111: c <= 9'b101001111;
				8'b101011: c <= 9'b10100;
				8'b1101011: c <= 9'b11111000;
				8'b111100: c <= 9'b1001011;
				8'b1000111: c <= 9'b1000110;
				8'b1011111: c <= 9'b10111011;
				8'b1110100: c <= 9'b101110010;
				8'b101101: c <= 9'b1101010;
				8'b1010011: c <= 9'b111100001;
				8'b1100001: c <= 9'b110001000;
				8'b110101: c <= 9'b11010011;
				8'b1000100: c <= 9'b10101;
				8'b1010001: c <= 9'b11100110;
				8'b1010100: c <= 9'b100001111;
				8'b1100110: c <= 9'b1;
				8'b101010: c <= 9'b1111001;
				8'b1011110: c <= 9'b111011011;
				8'b1100111: c <= 9'b1000;
				8'b1011010: c <= 9'b11001010;
				8'b1000010: c <= 9'b1100111;
				8'b111101: c <= 9'b101001110;
				8'b110000: c <= 9'b1100001;
				8'b111110: c <= 9'b11001101;
				8'b1100010: c <= 9'b101111010;
				8'b1110000: c <= 9'b1110111;
				8'b1101001: c <= 9'b111000110;
				8'b1110011: c <= 9'b111101101;
				8'b1001100: c <= 9'b10100;
				8'b100001: c <= 9'b1111101;
				8'b1000110: c <= 9'b110110111;
				8'b1110010: c <= 9'b101001000;
				8'b1010000: c <= 9'b110111000;
				8'b1111010: c <= 9'b110110111;
				8'b1010101: c <= 9'b101101100;
				8'b111011: c <= 9'b10101110;
				8'b1001101: c <= 9'b101001110;
				8'b111111: c <= 9'b101101000;
				8'b1101110: c <= 9'b11100010;
				8'b1111011: c <= 9'b101010110;
				8'b1001011: c <= 9'b100011100;
				8'b1101111: c <= 9'b1101010;
				8'b1101000: c <= 9'b111000010;
				8'b101100: c <= 9'b110;
				8'b100100: c <= 9'b110011011;
				8'b1111000: c <= 9'b11111101;
				8'b1000101: c <= 9'b110111;
				8'b1011001: c <= 9'b111100101;
				8'b110100: c <= 9'b111111110;
				8'b1111001: c <= 9'b100011010;
				8'b1110001: c <= 9'b111001;
				8'b1001111: c <= 9'b110100111;
				8'b1100101: c <= 9'b110011011;
				8'b1111110: c <= 9'b11110110;
				8'b1111100: c <= 9'b11001000;
				8'b1010110: c <= 9'b10111101;
				8'b110010: c <= 9'b101010;
				8'b1101101: c <= 9'b1111111;
				8'b100011: c <= 9'b10000010;
				8'b1110101: c <= 9'b10111000;
				8'b1111101: c <= 9'b100;
				8'b101001: c <= 9'b101001100;
				8'b1010010: c <= 9'b110010101;
				8'b1011000: c <= 9'b1001;
				8'b101110: c <= 9'b11001111;
				8'b1000001: c <= 9'b100010101;
				default: c <= 9'b0;
			endcase

		endcase
	end
endmodule

